///*****************************************************
//Title:    sb_ice_syn.v library verilog models
//Design:   sb_ice_syn.v
//Author:  
//Function: Verilog behavioral models for 
//          sb_ice_syn.v synthesis library
//Company:  SiliconBlue Technologies, Inc.
//******************************************************
`timescale 1ps/1ps
module SB_CARRY (CO, I0, I1, CI);
input I0, I1, CI;
output CO;
reg CI_int;

   assign CO = (CI_int * I0) | (CI_int * I1) | (I0 * I1);

   always @(CI)
	if ((CI == 1'b0) || (CI == 1'b1))
		CI_int = CI;
	else
		CI_int = 1'b0; // take care of CI is not connected if the CI is an output from LUT instead of from another CARRY

`ifdef TIMINGCHECK
specify
   (CI *> CO) = (1.0, 1.0);   
   (I0 *> CO) = (1.0, 1.0);
   (I1 *> CO) = (1.0, 1.0);   
endspecify
`endif

endmodule
`timescale 1ps/1ps
module SB_CARRY_IN_MUX (carry_init_out, carry_init_in);
   parameter C_INIT = 2'b00;  //c[1:0]
output carry_init_out;
input carry_init_in;
wire [1:0] select_bits;
reg carry_init_out;
assign select_bits = {C_INIT};
   always @ (select_bits or carry_init_in)
      case (select_bits)
         2'b00 :  carry_init_out = 1'b0;
         2'b01 :  carry_init_out = 1'b1;
         2'b10 :  carry_init_out = carry_init_in;
//         2'b11 :  carry_init_out = carry_init_in;
         default  : carry_init_out = 1'b0;
      endcase

`ifdef TIMINGCHECK
specify
   (carry_init_in *> carry_init_out) = (1.0, 1.0);

endspecify
`endif
endmodule
`timescale 1ps/1ps
module SB_LUT4 (O, I0, I1, I2, I3);
   parameter LUT_INIT = 16'h0000;
input I0, I1, I2, I3;
output O;
wire [15:0] mask;

reg luts;
reg I3_in, I2_in, I1_in, I0_in;
initial
begin
  luts = 1'b0;
  I3_in = 1'b0;
  I2_in = 1'b0;
  I1_in = 1'b0;
  I0_in = 1'b0;
end
always @ (I3 or I2 or I1 or I0)
  begin
    I3_in = I3;
    I2_in = I2;
    I1_in = I1;
    I0_in = I0;
  end
assign mask = LUT_INIT;
assign O = luts;

reg tmp;
always @(I3_in or I2_in or I1_in or I0_in ) begin
   tmp = I3_in ^ I2_in ^ I1_in ^ I0_in;
   #0.01;
   if (tmp === 0 || tmp === 1)
      luts = mask[{I3_in, I2_in, I1_in, I0_in}];
   else
      luts = lut_mux ({lut_mux (mask[15:12], {I1_in, I0_in}), lut_mux (mask[11:8], {I1_in, I0_in}), lut_mux (mask[7:4], {I1_in, I0_in}), lut_mux (mask[3:0], {I1_in, I0_in})}, {I3_in, I2_in});
end

function lut_mux;
input [3:0] d;
input [1:0] s;
   begin
      if ((s[1]^s[0] ==1) || (s[1]^s[0] ==0))
         lut_mux = d[s];
      else if ((d[0] ^ d[1]) == 0 && (d[2] ^ d[3]) == 0 && (d[0] ^ d[2]) == 0)
         lut_mux = d[0];
      else if ((s[1] == 0) && (d[0] == d[1]))
         lut_mux = d[0];
      else if ((s[1] == 1) && (d[2] == d[3]))
         lut_mux = d[2];
      else if ((s[0] == 0) && (d[0] == d[2]))
         lut_mux = d[0];
      else if ((s[0] == 1) && (d[1] == d[3]))
         lut_mux = d[1];
      else
         lut_mux = 1'bx;
   end
endfunction

endmodule
`timescale 1ps/1ps
module SB_DFF (Q, C, D);
input D, C;
output Q;
reg Q = 0;
   always @(posedge C)
         Q <= D;
endmodule
`timescale 1ps/1ps
module SB_DFFSR (Q, C, D, R);
input D, R, C;
output Q;
reg Q = 0;
   always @(posedge C)
         if (R) Q <= 1'b0; else Q <= D;
endmodule
`timescale 1ps/1ps
module SB_DFFSS (Q, C, D, S);
input D, S, C;
output Q;
reg Q = 0;
   always @(posedge C)
         if (S) Q <= 1'b1; else Q <= D;
endmodule
`timescale 1ps/1ps
module SB_DFFR (Q, C, D, R);
input C, D, R;
output Q;
reg Q = 0;
   always @(posedge C or posedge R)
      if (R) Q <= 1'b0;
      else  Q <= D;
endmodule
`timescale 1ps/1ps
module SB_DFFS (Q, C, D, S);
input D, S, C;
output Q;
reg Q = 0;
   always @(posedge C or posedge S)
      if (S) Q <= 1'b1;
      else Q <= D;
endmodule
`timescale 1ps/1ps
module SB_DFFE (Q, C, E, D);
input D, C, E;
output Q;
assign (weak0, weak1) E =1'b1 ;
reg Q = 0;
   always @(posedge C)
         if (E) Q <= D;
endmodule
`timescale 1ps/1ps
module SB_DFFESR (Q, C, E, D, R);
input D, R, C, E;
output Q;
assign (weak0, weak1) E =1'b1 ;
reg Q = 0;
   always @(posedge C)
         if (E) 
            if (R) Q <= 1'b0; else Q <= D;
endmodule
`timescale 1ps/1ps
module SB_DFFESS (Q, C, E, D, S);
input D, S, C, E;
output Q;
assign (weak0, weak1) E =1'b1 ;
reg Q = 0;
   always @(posedge C)
         if (E) 
            if (S) Q <= 1'b1; else Q <= D;
endmodule
`timescale 1ps/1ps
module SB_DFFER (Q, C, E, D, R);
input C, D, R, E;
output Q;
assign (weak0, weak1) E =1'b1 ;
reg Q = 0;
   always @(posedge C or posedge R)
      if (R) Q <= 1'b0;
      else if (E) Q <= D;
endmodule
`timescale 1ps/1ps
module SB_DFFES (Q, C, E, D, S);
input D, S, C, E;
output Q;
assign (weak0, weak1) E =1'b1 ;
reg Q = 0;
   always @(posedge C or posedge S)
      if (S) Q <= 1'b1;
      else if (E) Q <= D;
endmodule
`timescale 1ps/1ps
module SB_DFFN (Q, C, D);
input D, C;
output Q;
reg Q = 0;
   always @(negedge C)
         Q <= D;
endmodule
`timescale 1ps/1ps
module SB_DFFNSR (Q, C, D, R);
input D, R, C;
output Q;
reg Q = 0;
   always @(negedge C)
         if (R) Q <= 1'b0; else Q <= D;
endmodule
`timescale 1ps/1ps
module SB_DFFNSS (Q, C, D, S);
input D, S, C;
output Q;
reg Q = 0;
   always @(negedge C)
         if (S) Q <= 1'b1; else Q <= D;
endmodule
`timescale 1ps/1ps
module SB_DFFNR (Q, C, D, R);
input C, D, R;
output Q;
reg Q = 0;
   always @(negedge C or posedge R)
      if (R) Q <= 1'b0;
      else  Q <= D;
endmodule
`timescale 1ps/1ps
module SB_DFFNS (Q, C, D, S);
input D, S, C;
output Q;
reg Q = 0;
   always @(negedge  C or posedge S)
      if (S) Q <= 1'b1;
      else Q <= D;
endmodule
`timescale 1ps/1ps
module SB_DFFNE (Q, C, E, D);
input D, C, E;
output Q;
assign (weak0, weak1) E =1'b1 ;
reg Q = 0;
   always @(negedge C)
         if (E) Q <= D;
endmodule
`timescale 1ps/1ps
module SB_DFFNESR (Q, C, E, D, R);
input D, R, C, E;
output Q;
assign (weak0, weak1) E =1'b1 ;
reg Q = 0;
   always @(negedge C)
         if (E) 
            if (R) Q <= 1'b0; else Q <= D;
endmodule
`timescale 1ps/1ps
module SB_DFFNESS (Q, C, E, D, S);
input D, S, C, E;
output Q;
assign (weak0, weak1) E =1'b1 ;
reg Q = 0;
   always @(negedge C)
         if (E) 
            if (S) Q <= 1'b1; else Q <= D;
endmodule
`timescale 1ps/1ps
module SB_DFFNER (Q, C, E, D, R);
input C, D, R, E;
output Q;
assign (weak0, weak1) E =1'b1 ;
reg Q = 0;
   always @(negedge C or posedge R)
      if (R) Q <= 1'b0;
      else if (E) Q <= D;
endmodule
`timescale 1ps/1ps
module SB_DFFNES (Q, C, E, D, S);
input D, S, C, E;
output Q;
assign (weak0, weak1) E =1'b1 ;
reg Q = 0;
   always @(negedge C or posedge S)
      if (S) Q <= 1'b1;
      else if (E) Q <= D;
endmodule

`timescale 1ps/1ps
module SB_RAM4KNR (RDATA, RCLKN, RCLKE, RE, RADDR, WCLK, WCLKE, WE, WADDR, MASK, WDATA);
output [15:0] RDATA;
input RCLKN;
input RCLKE;
input RE;
input [7:0] RADDR;
input WCLK;
input WCLKE;
input WE;
input [7:0] WADDR;
input [15:0] MASK;
input [15:0] WDATA;

parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

wire RCLK;
assign (weak0, weak1) RCLKE =1'b1 ;
assign (weak0, weak1) RE =1'b0 ;
assign (weak0, weak1) WCLKE =1'b1 ;
assign (weak0, weak1) WE =1'b0 ;
assign RCLK = ~RCLKN;

SB_RAM4K sb_ram4k_inst (
	.RDATA(RDATA),
	.RCLK(RCLK),
	.RCLKE(RCLKE),
	.RE(RE),
	.RADDR(RADDR),
	.WCLK(WCLK),
	.WCLKE(WCLKE),
	.WE(WE),
	.WADDR(WADDR),
	.MASK(MASK),
	.WDATA(WDATA));

defparam sb_ram4k_inst.INIT_0 = INIT_0;
defparam sb_ram4k_inst.INIT_1 = INIT_1;
defparam sb_ram4k_inst.INIT_2 = INIT_2;
defparam sb_ram4k_inst.INIT_3 = INIT_3;
defparam sb_ram4k_inst.INIT_4 = INIT_4;
defparam sb_ram4k_inst.INIT_5 = INIT_5;
defparam sb_ram4k_inst.INIT_6 = INIT_6;
defparam sb_ram4k_inst.INIT_7 = INIT_7;
defparam sb_ram4k_inst.INIT_8 = INIT_8;
defparam sb_ram4k_inst.INIT_9 = INIT_9;
defparam sb_ram4k_inst.INIT_A = INIT_A;
defparam sb_ram4k_inst.INIT_B = INIT_B;
defparam sb_ram4k_inst.INIT_C = INIT_C;
defparam sb_ram4k_inst.INIT_D = INIT_D;
defparam sb_ram4k_inst.INIT_E = INIT_E;
defparam sb_ram4k_inst.INIT_F = INIT_F;

`ifdef TIMINGCHECK
specify
   (RCLKN *> RDATA[0]) = (1.0, 1.0);
   (RCLKN *> RDATA[1]) = (1.0, 1.0);
   (RCLKN *> RDATA[2]) = (1.0, 1.0);
   (RCLKN *> RDATA[3]) = (1.0, 1.0);
   (RCLKN *> RDATA[4]) = (1.0, 1.0);
   (RCLKN *> RDATA[5]) = (1.0, 1.0);
   (RCLKN *> RDATA[6]) = (1.0, 1.0);
   (RCLKN *> RDATA[7]) = (1.0, 1.0);
   (RCLKN *> RDATA[8]) = (1.0, 1.0);
   (RCLKN *> RDATA[9]) = (1.0, 1.0);
   (RCLKN *> RDATA[10]) = (1.0, 1.0);
   (RCLKN *> RDATA[11]) = (1.0, 1.0);
   (RCLKN *> RDATA[12]) = (1.0, 1.0);
   (RCLKN *> RDATA[13]) = (1.0, 1.0);
   (RCLKN *> RDATA[14]) = (1.0, 1.0);
   (RCLKN *> RDATA[15]) = (1.0, 1.0);
   $setup(posedge MASK[0], posedge WCLK, 1.0);
   $setup(negedge MASK[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[0], 1.0);
   $hold(posedge WCLK, negedge MASK[0], 1.0);
   $setup(posedge MASK[1], posedge WCLK, 1.0);
   $setup(negedge MASK[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[1], 1.0);
   $hold(posedge WCLK, negedge MASK[1], 1.0);
   $setup(posedge MASK[2], posedge WCLK, 1.0);
   $setup(negedge MASK[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[2], 1.0);
   $hold(posedge WCLK, negedge MASK[2], 1.0);
   $setup(posedge MASK[3], posedge WCLK, 1.0);
   $setup(negedge MASK[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[3], 1.0);
   $hold(posedge WCLK, negedge MASK[3], 1.0);
   $setup(posedge MASK[4], posedge WCLK, 1.0);
   $setup(negedge MASK[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[4], 1.0);
   $hold(posedge WCLK, negedge MASK[4], 1.0);
   $setup(posedge MASK[5], posedge WCLK, 1.0);
   $setup(negedge MASK[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[5], 1.0);
   $hold(posedge WCLK, negedge MASK[5], 1.0);
   $setup(posedge MASK[6], posedge WCLK, 1.0);
   $setup(negedge MASK[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[6], 1.0);
   $hold(posedge WCLK, negedge MASK[6], 1.0);
   $setup(posedge MASK[7], posedge WCLK, 1.0);
   $setup(negedge MASK[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[7], 1.0);
   $hold(posedge WCLK, negedge MASK[7], 1.0);
   $setup(posedge MASK[8], posedge WCLK, 1.0);
   $setup(negedge MASK[8], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[8], 1.0);
   $hold(posedge WCLK, negedge MASK[8], 1.0);
   $setup(posedge MASK[9], posedge WCLK, 1.0);
   $setup(negedge MASK[9], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[9], 1.0);
   $hold(posedge WCLK, negedge MASK[9], 1.0);
   $setup(posedge MASK[10], posedge WCLK, 1.0);
   $setup(negedge MASK[10], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[10], 1.0);
   $hold(posedge WCLK, negedge MASK[10], 1.0);
   $setup(posedge MASK[11], posedge WCLK, 1.0);
   $setup(negedge MASK[11], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[11], 1.0);
   $hold(posedge WCLK, negedge MASK[11], 1.0);
   $setup(posedge MASK[12], posedge WCLK, 1.0);
   $setup(negedge MASK[12], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[12], 1.0);
   $hold(posedge WCLK, negedge MASK[12], 1.0);
   $setup(posedge MASK[13], posedge WCLK, 1.0);
   $setup(negedge MASK[13], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[13], 1.0);
   $hold(posedge WCLK, negedge MASK[13], 1.0);
   $setup(posedge MASK[14], posedge WCLK, 1.0);
   $setup(negedge MASK[14], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[14], 1.0);
   $hold(posedge WCLK, negedge MASK[14], 1.0);
   $setup(posedge MASK[15], posedge WCLK, 1.0);
   $setup(negedge MASK[15], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[15], 1.0);
   $hold(posedge WCLK, negedge MASK[15], 1.0);
   $setup(posedge WADDR[0], posedge WCLK, 1.0);
   $setup(negedge WADDR[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[0], 1.0);
   $hold(posedge WCLK, negedge WADDR[0], 1.0);
   $setup(posedge WADDR[1], posedge WCLK, 1.0);
   $setup(negedge WADDR[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[1], 1.0);
   $hold(posedge WCLK, negedge WADDR[1], 1.0);
   $setup(posedge WADDR[2], posedge WCLK, 1.0);
   $setup(negedge WADDR[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[2], 1.0);
   $hold(posedge WCLK, negedge WADDR[2], 1.0);
   $setup(posedge WADDR[3], posedge WCLK, 1.0);
   $setup(negedge WADDR[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[3], 1.0);
   $hold(posedge WCLK, negedge WADDR[3], 1.0);
   $setup(posedge WADDR[4], posedge WCLK, 1.0);
   $setup(negedge WADDR[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[4], 1.0);
   $hold(posedge WCLK, negedge WADDR[4], 1.0);
   $setup(posedge WADDR[5], posedge WCLK, 1.0);
   $setup(negedge WADDR[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[5], 1.0);
   $hold(posedge WCLK, negedge WADDR[5], 1.0);
   $setup(posedge WADDR[6], posedge WCLK, 1.0);
   $setup(negedge WADDR[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[6], 1.0);
   $hold(posedge WCLK, negedge WADDR[6], 1.0);
   $setup(posedge WADDR[7], posedge WCLK, 1.0);
   $setup(negedge WADDR[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[7], 1.0);
   $hold(posedge WCLK, negedge WADDR[7], 1.0);
   $setup(posedge WDATA[0], posedge WCLK, 1.0);
   $setup(negedge WDATA[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[0], 1.0);
   $hold(posedge WCLK, negedge WDATA[0], 1.0);
   $setup(posedge WDATA[1], posedge WCLK, 1.0);
   $setup(negedge WDATA[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[1], 1.0);
   $hold(posedge WCLK, negedge WDATA[1], 1.0);
   $setup(posedge WDATA[2], posedge WCLK, 1.0);
   $setup(negedge WDATA[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[2], 1.0);
   $hold(posedge WCLK, negedge WDATA[2], 1.0);
   $setup(posedge WDATA[3], posedge WCLK, 1.0);
   $setup(negedge WDATA[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[3], 1.0);
   $hold(posedge WCLK, negedge WDATA[3], 1.0);
   $setup(posedge WDATA[4], posedge WCLK, 1.0);
   $setup(negedge WDATA[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[4], 1.0);
   $hold(posedge WCLK, negedge WDATA[4], 1.0);
   $setup(posedge WDATA[5], posedge WCLK, 1.0);
   $setup(negedge WDATA[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[5], 1.0);
   $hold(posedge WCLK, negedge WDATA[5], 1.0);
   $setup(posedge WDATA[6], posedge WCLK, 1.0);
   $setup(negedge WDATA[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[6], 1.0);
   $hold(posedge WCLK, negedge WDATA[6], 1.0);
   $setup(posedge WDATA[7], posedge WCLK, 1.0);
   $setup(negedge WDATA[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[7], 1.0);
   $hold(posedge WCLK, negedge WDATA[7], 1.0);
   $setup(posedge WDATA[8], posedge WCLK, 1.0);
   $setup(negedge WDATA[8], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[8], 1.0);
   $hold(posedge WCLK, negedge WDATA[8], 1.0);
   $setup(posedge WDATA[9], posedge WCLK, 1.0);
   $setup(negedge WDATA[9], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[9], 1.0);
   $hold(posedge WCLK, negedge WDATA[9], 1.0);
   $setup(posedge WDATA[10], posedge WCLK, 1.0);
   $setup(negedge WDATA[10], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[10], 1.0);
   $hold(posedge WCLK, negedge WDATA[10], 1.0);
   $setup(posedge WDATA[11], posedge WCLK, 1.0);
   $setup(negedge WDATA[11], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[11], 1.0);
   $hold(posedge WCLK, negedge WDATA[11], 1.0);
   $setup(posedge WDATA[12], posedge WCLK, 1.0);
   $setup(negedge WDATA[12], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[12], 1.0);
   $hold(posedge WCLK, negedge WDATA[12], 1.0);
   $setup(posedge WDATA[13], posedge WCLK, 1.0);
   $setup(negedge WDATA[13], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[13], 1.0);
   $hold(posedge WCLK, negedge WDATA[13], 1.0);
   $setup(posedge WDATA[14], posedge WCLK, 1.0);
   $setup(negedge WDATA[14], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[14], 1.0);
   $hold(posedge WCLK, negedge WDATA[14], 1.0);
   $setup(posedge WDATA[15], posedge WCLK, 1.0);
   $setup(negedge WDATA[15], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[15], 1.0);
   $hold(posedge WCLK, negedge WDATA[15], 1.0);
   $setup(posedge WCLKE, posedge WCLK, 1.0);
   $setup(negedge WCLKE, posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WCLKE, 1.0);
   $hold(posedge WCLK, negedge WCLKE, 1.0);
   $setup(posedge WE, posedge WCLK, 1.0);
   $setup(negedge WE, posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WE, 1.0);
   $hold(posedge WCLK, negedge WE, 1.0);
   $setup(posedge RADDR[0], posedge RCLKN, 1.0);
   $setup(negedge RADDR[0], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[0], 1.0);
   $hold(posedge RCLKN, negedge RADDR[0], 1.0);
   $setup(posedge RADDR[1], posedge RCLKN, 1.0);
   $setup(negedge RADDR[1], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[1], 1.0);
   $hold(posedge RCLKN, negedge RADDR[1], 1.0);
   $setup(posedge RADDR[2], posedge RCLKN, 1.0);
   $setup(negedge RADDR[2], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[2], 1.0);
   $hold(posedge RCLKN, negedge RADDR[2], 1.0);
   $setup(posedge RADDR[3], posedge RCLKN, 1.0);
   $setup(negedge RADDR[3], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[3], 1.0);
   $hold(posedge RCLKN, negedge RADDR[3], 1.0);
   $setup(posedge RADDR[4], posedge RCLKN, 1.0);
   $setup(negedge RADDR[4], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[4], 1.0);
   $hold(posedge RCLKN, negedge RADDR[4], 1.0);
   $setup(posedge RADDR[5], posedge RCLKN, 1.0);
   $setup(negedge RADDR[5], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[5], 1.0);
   $hold(posedge RCLKN, negedge RADDR[5], 1.0);
   $setup(posedge RADDR[6], posedge RCLKN, 1.0);
   $setup(negedge RADDR[6], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[6], 1.0);
   $hold(posedge RCLKN, negedge RADDR[6], 1.0);
   $setup(posedge RADDR[7], posedge RCLKN, 1.0);
   $setup(negedge RADDR[7], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[7], 1.0);
   $hold(posedge RCLKN, negedge RADDR[7], 1.0);
   $setup(posedge RCLKE, posedge RCLKN, 1.0);
   $setup(negedge RCLKE, posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RCLKE, 1.0);
   $hold(posedge RCLKN, negedge RCLKE, 1.0);
   $setup(posedge RE, posedge RCLKN, 1.0);
   $setup(negedge RE, posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RE, 1.0);
   $hold(posedge RCLKN, negedge RE, 1.0);
   $recovery(posedge RCLKN, posedge WCLK, 1.0);
   $recovery(negedge RCLKN, posedge WCLK, 1.0);
   $removal(posedge RCLKN, posedge WCLK, 1.0);
   $removal(negedge RCLKN, posedge WCLK, 1.0);
   $recovery(posedge WCLK, posedge RCLKN, 1.0);
   $recovery(negedge WCLK, posedge RCLKN, 1.0);
   $removal(posedge WCLK, posedge RCLKN, 1.0);
   $removal(negedge WCLK, posedge RCLKN, 1.0);

endspecify
`endif

endmodule //SB_RAM4KNR
`timescale 1ps/1ps
module SB_RAM4KNW (RDATA, RCLK, RCLKE, RE, RADDR, WCLKN, WCLKE, WE, WADDR, MASK, WDATA);
output [15:0] RDATA;
input RCLK;
input RCLKE;
input RE;
input [7:0] RADDR;
input WCLKN;
input WCLKE;
input WE;
input [7:0] WADDR;
input [15:0] MASK;
input [15:0] WDATA;

parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

wire WCLK;
assign (weak0, weak1) RCLKE =1'b1 ;
assign (weak0, weak1) RE =1'b0 ;
assign (weak0, weak1) WCLKE =1'b1 ;
assign (weak0, weak1) WE =1'b0 ;
assign WCLK = ~WCLKN;

SB_RAM4K sb_ram4k_inst (
	.RDATA(RDATA),
	.RCLK(RCLK),
	.RCLKE(RCLKE),
	.RE(RE),
	.RADDR(RADDR),
	.WCLK(WCLK),
	.WCLKE(WCLKE),
	.WE(WE),
	.WADDR(WADDR),
	.MASK(MASK),
	.WDATA(WDATA));

defparam sb_ram4k_inst.INIT_0 = INIT_0;
defparam sb_ram4k_inst.INIT_1 = INIT_1;
defparam sb_ram4k_inst.INIT_2 = INIT_2;
defparam sb_ram4k_inst.INIT_3 = INIT_3;
defparam sb_ram4k_inst.INIT_4 = INIT_4;
defparam sb_ram4k_inst.INIT_5 = INIT_5;
defparam sb_ram4k_inst.INIT_6 = INIT_6;
defparam sb_ram4k_inst.INIT_7 = INIT_7;
defparam sb_ram4k_inst.INIT_8 = INIT_8;
defparam sb_ram4k_inst.INIT_9 = INIT_9;
defparam sb_ram4k_inst.INIT_A = INIT_A;
defparam sb_ram4k_inst.INIT_B = INIT_B;
defparam sb_ram4k_inst.INIT_C = INIT_C;
defparam sb_ram4k_inst.INIT_D = INIT_D;
defparam sb_ram4k_inst.INIT_E = INIT_E;
defparam sb_ram4k_inst.INIT_F = INIT_F;

`ifdef TIMINGCHECK
specify
   (RCLK *> RDATA[0]) = (1.0, 1.0);
   (RCLK *> RDATA[1]) = (1.0, 1.0);
   (RCLK *> RDATA[2]) = (1.0, 1.0);
   (RCLK *> RDATA[3]) = (1.0, 1.0);
   (RCLK *> RDATA[4]) = (1.0, 1.0);
   (RCLK *> RDATA[5]) = (1.0, 1.0);
   (RCLK *> RDATA[6]) = (1.0, 1.0);
   (RCLK *> RDATA[7]) = (1.0, 1.0);
   (RCLK *> RDATA[8]) = (1.0, 1.0);
   (RCLK *> RDATA[9]) = (1.0, 1.0);
   (RCLK *> RDATA[10]) = (1.0, 1.0);
   (RCLK *> RDATA[11]) = (1.0, 1.0);
   (RCLK *> RDATA[12]) = (1.0, 1.0);
   (RCLK *> RDATA[13]) = (1.0, 1.0);
   (RCLK *> RDATA[14]) = (1.0, 1.0);
   (RCLK *> RDATA[15]) = (1.0, 1.0);
   $setup(posedge MASK[0], posedge WCLKN, 1.0);
   $setup(negedge MASK[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[0], 1.0);
   $hold(posedge WCLKN, negedge MASK[0], 1.0);
   $setup(posedge MASK[1], posedge WCLKN, 1.0);
   $setup(negedge MASK[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[1], 1.0);
   $hold(posedge WCLKN, negedge MASK[1], 1.0);
   $setup(posedge MASK[2], posedge WCLKN, 1.0);
   $setup(negedge MASK[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[2], 1.0);
   $hold(posedge WCLKN, negedge MASK[2], 1.0);
   $setup(posedge MASK[3], posedge WCLKN, 1.0);
   $setup(negedge MASK[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[3], 1.0);
   $hold(posedge WCLKN, negedge MASK[3], 1.0);
   $setup(posedge MASK[4], posedge WCLKN, 1.0);
   $setup(negedge MASK[4], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[4], 1.0);
   $hold(posedge WCLKN, negedge MASK[4], 1.0);
   $setup(posedge MASK[5], posedge WCLKN, 1.0);
   $setup(negedge MASK[5], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[5], 1.0);
   $hold(posedge WCLKN, negedge MASK[5], 1.0);
   $setup(posedge MASK[6], posedge WCLKN, 1.0);
   $setup(negedge MASK[6], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[6], 1.0);
   $hold(posedge WCLKN, negedge MASK[6], 1.0);
   $setup(posedge MASK[7], posedge WCLKN, 1.0);
   $setup(negedge MASK[7], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[7], 1.0);
   $hold(posedge WCLKN, negedge MASK[7], 1.0);
   $setup(posedge MASK[8], posedge WCLKN, 1.0);
   $setup(negedge MASK[8], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[8], 1.0);
   $hold(posedge WCLKN, negedge MASK[8], 1.0);
   $setup(posedge MASK[9], posedge WCLKN, 1.0);
   $setup(negedge MASK[9], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[9], 1.0);
   $hold(posedge WCLKN, negedge MASK[9], 1.0);
   $setup(posedge MASK[10], posedge WCLKN, 1.0);
   $setup(negedge MASK[10], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[10], 1.0);
   $hold(posedge WCLKN, negedge MASK[10], 1.0);
   $setup(posedge MASK[11], posedge WCLKN, 1.0);
   $setup(negedge MASK[11], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[11], 1.0);
   $hold(posedge WCLKN, negedge MASK[11], 1.0);
   $setup(posedge MASK[12], posedge WCLKN, 1.0);
   $setup(negedge MASK[12], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[12], 1.0);
   $hold(posedge WCLKN, negedge MASK[12], 1.0);
   $setup(posedge MASK[13], posedge WCLKN, 1.0);
   $setup(negedge MASK[13], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[13], 1.0);
   $hold(posedge WCLKN, negedge MASK[13], 1.0);
   $setup(posedge MASK[14], posedge WCLKN, 1.0);
   $setup(negedge MASK[14], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[14], 1.0);
   $hold(posedge WCLKN, negedge MASK[14], 1.0);
   $setup(posedge MASK[15], posedge WCLKN, 1.0);
   $setup(negedge MASK[15], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[15], 1.0);
   $hold(posedge WCLKN, negedge MASK[15], 1.0);
   $setup(posedge WADDR[0], posedge WCLKN, 1.0);
   $setup(negedge WADDR[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[0], 1.0);
   $hold(posedge WCLKN, negedge WADDR[0], 1.0);
   $setup(posedge WADDR[1], posedge WCLKN, 1.0);
   $setup(negedge WADDR[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[1], 1.0);
   $hold(posedge WCLKN, negedge WADDR[1], 1.0);
   $setup(posedge WADDR[2], posedge WCLKN, 1.0);
   $setup(negedge WADDR[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[2], 1.0);
   $hold(posedge WCLKN, negedge WADDR[2], 1.0);
   $setup(posedge WADDR[3], posedge WCLKN, 1.0);
   $setup(negedge WADDR[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[3], 1.0);
   $hold(posedge WCLKN, negedge WADDR[3], 1.0);
   $setup(posedge WADDR[4], posedge WCLKN, 1.0);
   $setup(negedge WADDR[4], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[4], 1.0);
   $hold(posedge WCLKN, negedge WADDR[4], 1.0);
   $setup(posedge WADDR[5], posedge WCLKN, 1.0);
   $setup(negedge WADDR[5], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[5], 1.0);
   $hold(posedge WCLKN, negedge WADDR[5], 1.0);
   $setup(posedge WADDR[6], posedge WCLKN, 1.0);
   $setup(negedge WADDR[6], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[6], 1.0);
   $hold(posedge WCLKN, negedge WADDR[6], 1.0);
   $setup(posedge WADDR[7], posedge WCLKN, 1.0);
   $setup(negedge WADDR[7], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[7], 1.0);
   $hold(posedge WCLKN, negedge WADDR[7], 1.0);
   $setup(posedge WDATA[0], posedge WCLKN, 1.0);
   $setup(negedge WDATA[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[0], 1.0);
   $hold(posedge WCLKN, negedge WDATA[0], 1.0);
   $setup(posedge WDATA[1], posedge WCLKN, 1.0);
   $setup(negedge WDATA[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[1], 1.0);
   $hold(posedge WCLKN, negedge WDATA[1], 1.0);
   $setup(posedge WDATA[2], posedge WCLKN, 1.0);
   $setup(negedge WDATA[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[2], 1.0);
   $hold(posedge WCLKN, negedge WDATA[2], 1.0);
   $setup(posedge WDATA[3], posedge WCLKN, 1.0);
   $setup(negedge WDATA[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[3], 1.0);
   $hold(posedge WCLKN, negedge WDATA[3], 1.0);
   $setup(posedge WDATA[4], posedge WCLKN, 1.0);
   $setup(negedge WDATA[4], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[4], 1.0);
   $hold(posedge WCLKN, negedge WDATA[4], 1.0);
   $setup(posedge WDATA[5], posedge WCLKN, 1.0);
   $setup(negedge WDATA[5], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[5], 1.0);
   $hold(posedge WCLKN, negedge WDATA[5], 1.0);
   $setup(posedge WDATA[6], posedge WCLKN, 1.0);
   $setup(negedge WDATA[6], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[6], 1.0);
   $hold(posedge WCLKN, negedge WDATA[6], 1.0);
   $setup(posedge WDATA[7], posedge WCLKN, 1.0);
   $setup(negedge WDATA[7], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[7], 1.0);
   $hold(posedge WCLKN, negedge WDATA[7], 1.0);
   $setup(posedge WDATA[8], posedge WCLKN, 1.0);
   $setup(negedge WDATA[8], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[8], 1.0);
   $hold(posedge WCLKN, negedge WDATA[8], 1.0);
   $setup(posedge WDATA[9], posedge WCLKN, 1.0);
   $setup(negedge WDATA[9], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[9], 1.0);
   $hold(posedge WCLKN, negedge WDATA[9], 1.0);
   $setup(posedge WDATA[10], posedge WCLKN, 1.0);
   $setup(negedge WDATA[10], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[10], 1.0);
   $hold(posedge WCLKN, negedge WDATA[10], 1.0);
   $setup(posedge WDATA[11], posedge WCLKN, 1.0);
   $setup(negedge WDATA[11], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[11], 1.0);
   $hold(posedge WCLKN, negedge WDATA[11], 1.0);
   $setup(posedge WDATA[12], posedge WCLKN, 1.0);
   $setup(negedge WDATA[12], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[12], 1.0);
   $hold(posedge WCLKN, negedge WDATA[12], 1.0);
   $setup(posedge WDATA[13], posedge WCLKN, 1.0);
   $setup(negedge WDATA[13], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[13], 1.0);
   $hold(posedge WCLKN, negedge WDATA[13], 1.0);
   $setup(posedge WDATA[14], posedge WCLKN, 1.0);
   $setup(negedge WDATA[14], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[14], 1.0);
   $hold(posedge WCLKN, negedge WDATA[14], 1.0);
   $setup(posedge WDATA[15], posedge WCLKN, 1.0);
   $setup(negedge WDATA[15], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[15], 1.0);
   $hold(posedge WCLKN, negedge WDATA[15], 1.0);
   $setup(posedge WCLKE, posedge WCLKN, 1.0);
   $setup(negedge WCLKE, posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WCLKE, 1.0);
   $hold(posedge WCLKN, negedge WCLKE, 1.0);
   $setup(posedge WE, posedge WCLKN, 1.0);
   $setup(negedge WE, posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WE, 1.0);
   $hold(posedge WCLKN, negedge WE, 1.0);
   $setup(posedge RADDR[0], posedge RCLK, 1.0);
   $setup(negedge RADDR[0], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[0], 1.0);
   $hold(posedge RCLK, negedge RADDR[0], 1.0);
   $setup(posedge RADDR[1], posedge RCLK, 1.0);
   $setup(negedge RADDR[1], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[1], 1.0);
   $hold(posedge RCLK, negedge RADDR[1], 1.0);
   $setup(posedge RADDR[2], posedge RCLK, 1.0);
   $setup(negedge RADDR[2], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[2], 1.0);
   $hold(posedge RCLK, negedge RADDR[2], 1.0);
   $setup(posedge RADDR[3], posedge RCLK, 1.0);
   $setup(negedge RADDR[3], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[3], 1.0);
   $hold(posedge RCLK, negedge RADDR[3], 1.0);
   $setup(posedge RADDR[4], posedge RCLK, 1.0);
   $setup(negedge RADDR[4], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[4], 1.0);
   $hold(posedge RCLK, negedge RADDR[4], 1.0);
   $setup(posedge RADDR[5], posedge RCLK, 1.0);
   $setup(negedge RADDR[5], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[5], 1.0);
   $hold(posedge RCLK, negedge RADDR[5], 1.0);
   $setup(posedge RADDR[6], posedge RCLK, 1.0);
   $setup(negedge RADDR[6], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[6], 1.0);
   $hold(posedge RCLK, negedge RADDR[6], 1.0);
   $setup(posedge RADDR[7], posedge RCLK, 1.0);
   $setup(negedge RADDR[7], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[7], 1.0);
   $hold(posedge RCLK, negedge RADDR[7], 1.0);
   $setup(posedge RCLKE, posedge RCLK, 1.0);
   $setup(negedge RCLKE, posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RCLKE, 1.0);
   $hold(posedge RCLK, negedge RCLKE, 1.0);
   $setup(posedge RE, posedge RCLK, 1.0);
   $setup(negedge RE, posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RE, 1.0);
   $hold(posedge RCLK, negedge RE, 1.0);
   $recovery(posedge RCLK, posedge WCLKN, 1.0);
   $recovery(negedge RCLK, posedge WCLKN, 1.0);
   $removal(posedge RCLK, posedge WCLKN, 1.0);
   $removal(negedge RCLK, posedge WCLKN, 1.0);
   $recovery(posedge WCLKN, posedge RCLK, 1.0);
   $recovery(negedge WCLKN, posedge RCLK, 1.0);
   $removal(posedge WCLKN, posedge RCLK, 1.0);
   $removal(negedge WCLKN, posedge RCLK, 1.0);

endspecify
`endif

endmodule //SB_RAM4KNW
`timescale 1ps/1ps
module SB_RAM4KNRNW (RDATA, RCLKN, RCLKE, RE, RADDR, WCLKN, WCLKE, WE, WADDR, MASK, WDATA);
output [15:0] RDATA;
input RCLKN;
input RCLKE;
input RE;
input [7:0] RADDR;
input WCLKN;
input WCLKE;
input WE;
input [7:0] WADDR;
input [15:0] MASK;
input [15:0] WDATA;

parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

wire RCLK, WCLK;
assign (weak0, weak1) RCLKE =1'b1 ;
assign (weak0, weak1) RE =1'b0 ;
assign (weak0, weak1) WCLKE =1'b1 ;
assign (weak0, weak1) WE =1'b0 ;
assign RCLK = ~RCLKN;
assign WCLK = ~WCLKN;

SB_RAM4K sb_ram4k_inst (
	.RDATA(RDATA),
	.RCLK(RCLK),
	.RCLKE(RCLKE),
	.RE(RE),
	.RADDR(RADDR),
	.WCLK(WCLK),
	.WCLKE(WCLKE),
	.WE(WE),
	.WADDR(WADDR),
	.MASK(MASK),
	.WDATA(WDATA));

defparam sb_ram4k_inst.INIT_0 = INIT_0;
defparam sb_ram4k_inst.INIT_1 = INIT_1;
defparam sb_ram4k_inst.INIT_2 = INIT_2;
defparam sb_ram4k_inst.INIT_3 = INIT_3;
defparam sb_ram4k_inst.INIT_4 = INIT_4;
defparam sb_ram4k_inst.INIT_5 = INIT_5;
defparam sb_ram4k_inst.INIT_6 = INIT_6;
defparam sb_ram4k_inst.INIT_7 = INIT_7;
defparam sb_ram4k_inst.INIT_8 = INIT_8;
defparam sb_ram4k_inst.INIT_9 = INIT_9;
defparam sb_ram4k_inst.INIT_A = INIT_A;
defparam sb_ram4k_inst.INIT_B = INIT_B;
defparam sb_ram4k_inst.INIT_C = INIT_C;
defparam sb_ram4k_inst.INIT_D = INIT_D;
defparam sb_ram4k_inst.INIT_E = INIT_E;
defparam sb_ram4k_inst.INIT_F = INIT_F;

`ifdef TIMINGCHECK
specify
   (RCLKN *> RDATA[0]) = (1.0, 1.0);
   (RCLKN *> RDATA[1]) = (1.0, 1.0);
   (RCLKN *> RDATA[2]) = (1.0, 1.0);
   (RCLKN *> RDATA[3]) = (1.0, 1.0);
   (RCLKN *> RDATA[4]) = (1.0, 1.0);
   (RCLKN *> RDATA[5]) = (1.0, 1.0);
   (RCLKN *> RDATA[6]) = (1.0, 1.0);
   (RCLKN *> RDATA[7]) = (1.0, 1.0);
   (RCLKN *> RDATA[8]) = (1.0, 1.0);
   (RCLKN *> RDATA[9]) = (1.0, 1.0);
   (RCLKN *> RDATA[10]) = (1.0, 1.0);
   (RCLKN *> RDATA[11]) = (1.0, 1.0);
   (RCLKN *> RDATA[12]) = (1.0, 1.0);
   (RCLKN *> RDATA[13]) = (1.0, 1.0);
   (RCLKN *> RDATA[14]) = (1.0, 1.0);
   (RCLKN *> RDATA[15]) = (1.0, 1.0);
   $setup(posedge MASK[0], posedge WCLKN, 1.0);
   $setup(negedge MASK[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[0], 1.0);
   $hold(posedge WCLKN, negedge MASK[0], 1.0);
   $setup(posedge MASK[1], posedge WCLKN, 1.0);
   $setup(negedge MASK[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[1], 1.0);
   $hold(posedge WCLKN, negedge MASK[1], 1.0);
   $setup(posedge MASK[2], posedge WCLKN, 1.0);
   $setup(negedge MASK[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[2], 1.0);
   $hold(posedge WCLKN, negedge MASK[2], 1.0);
   $setup(posedge MASK[3], posedge WCLKN, 1.0);
   $setup(negedge MASK[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[3], 1.0);
   $hold(posedge WCLKN, negedge MASK[3], 1.0);
   $setup(posedge MASK[4], posedge WCLKN, 1.0);
   $setup(negedge MASK[4], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[4], 1.0);
   $hold(posedge WCLKN, negedge MASK[4], 1.0);
   $setup(posedge MASK[5], posedge WCLKN, 1.0);
   $setup(negedge MASK[5], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[5], 1.0);
   $hold(posedge WCLKN, negedge MASK[5], 1.0);
   $setup(posedge MASK[6], posedge WCLKN, 1.0);
   $setup(negedge MASK[6], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[6], 1.0);
   $hold(posedge WCLKN, negedge MASK[6], 1.0);
   $setup(posedge MASK[7], posedge WCLKN, 1.0);
   $setup(negedge MASK[7], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[7], 1.0);
   $hold(posedge WCLKN, negedge MASK[7], 1.0);
   $setup(posedge MASK[8], posedge WCLKN, 1.0);
   $setup(negedge MASK[8], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[8], 1.0);
   $hold(posedge WCLKN, negedge MASK[8], 1.0);
   $setup(posedge MASK[9], posedge WCLKN, 1.0);
   $setup(negedge MASK[9], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[9], 1.0);
   $hold(posedge WCLKN, negedge MASK[9], 1.0);
   $setup(posedge MASK[10], posedge WCLKN, 1.0);
   $setup(negedge MASK[10], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[10], 1.0);
   $hold(posedge WCLKN, negedge MASK[10], 1.0);
   $setup(posedge MASK[11], posedge WCLKN, 1.0);
   $setup(negedge MASK[11], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[11], 1.0);
   $hold(posedge WCLKN, negedge MASK[11], 1.0);
   $setup(posedge MASK[12], posedge WCLKN, 1.0);
   $setup(negedge MASK[12], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[12], 1.0);
   $hold(posedge WCLKN, negedge MASK[12], 1.0);
   $setup(posedge MASK[13], posedge WCLKN, 1.0);
   $setup(negedge MASK[13], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[13], 1.0);
   $hold(posedge WCLKN, negedge MASK[13], 1.0);
   $setup(posedge MASK[14], posedge WCLKN, 1.0);
   $setup(negedge MASK[14], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[14], 1.0);
   $hold(posedge WCLKN, negedge MASK[14], 1.0);
   $setup(posedge MASK[15], posedge WCLKN, 1.0);
   $setup(negedge MASK[15], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[15], 1.0);
   $hold(posedge WCLKN, negedge MASK[15], 1.0);
   $setup(posedge WADDR[0], posedge WCLKN, 1.0);
   $setup(negedge WADDR[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[0], 1.0);
   $hold(posedge WCLKN, negedge WADDR[0], 1.0);
   $setup(posedge WADDR[1], posedge WCLKN, 1.0);
   $setup(negedge WADDR[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[1], 1.0);
   $hold(posedge WCLKN, negedge WADDR[1], 1.0);
   $setup(posedge WADDR[2], posedge WCLKN, 1.0);
   $setup(negedge WADDR[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[2], 1.0);
   $hold(posedge WCLKN, negedge WADDR[2], 1.0);
   $setup(posedge WADDR[3], posedge WCLKN, 1.0);
   $setup(negedge WADDR[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[3], 1.0);
   $hold(posedge WCLKN, negedge WADDR[3], 1.0);
   $setup(posedge WADDR[4], posedge WCLKN, 1.0);
   $setup(negedge WADDR[4], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[4], 1.0);
   $hold(posedge WCLKN, negedge WADDR[4], 1.0);
   $setup(posedge WADDR[5], posedge WCLKN, 1.0);
   $setup(negedge WADDR[5], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[5], 1.0);
   $hold(posedge WCLKN, negedge WADDR[5], 1.0);
   $setup(posedge WADDR[6], posedge WCLKN, 1.0);
   $setup(negedge WADDR[6], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[6], 1.0);
   $hold(posedge WCLKN, negedge WADDR[6], 1.0);
   $setup(posedge WADDR[7], posedge WCLKN, 1.0);
   $setup(negedge WADDR[7], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[7], 1.0);
   $hold(posedge WCLKN, negedge WADDR[7], 1.0);
   $setup(posedge WDATA[0], posedge WCLKN, 1.0);
   $setup(negedge WDATA[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[0], 1.0);
   $hold(posedge WCLKN, negedge WDATA[0], 1.0);
   $setup(posedge WDATA[1], posedge WCLKN, 1.0);
   $setup(negedge WDATA[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[1], 1.0);
   $hold(posedge WCLKN, negedge WDATA[1], 1.0);
   $setup(posedge WDATA[2], posedge WCLKN, 1.0);
   $setup(negedge WDATA[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[2], 1.0);
   $hold(posedge WCLKN, negedge WDATA[2], 1.0);
   $setup(posedge WDATA[3], posedge WCLKN, 1.0);
   $setup(negedge WDATA[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[3], 1.0);
   $hold(posedge WCLKN, negedge WDATA[3], 1.0);
   $setup(posedge WDATA[4], posedge WCLKN, 1.0);
   $setup(negedge WDATA[4], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[4], 1.0);
   $hold(posedge WCLKN, negedge WDATA[4], 1.0);
   $setup(posedge WDATA[5], posedge WCLKN, 1.0);
   $setup(negedge WDATA[5], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[5], 1.0);
   $hold(posedge WCLKN, negedge WDATA[5], 1.0);
   $setup(posedge WDATA[6], posedge WCLKN, 1.0);
   $setup(negedge WDATA[6], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[6], 1.0);
   $hold(posedge WCLKN, negedge WDATA[6], 1.0);
   $setup(posedge WDATA[7], posedge WCLKN, 1.0);
   $setup(negedge WDATA[7], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[7], 1.0);
   $hold(posedge WCLKN, negedge WDATA[7], 1.0);
   $setup(posedge WDATA[8], posedge WCLKN, 1.0);
   $setup(negedge WDATA[8], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[8], 1.0);
   $hold(posedge WCLKN, negedge WDATA[8], 1.0);
   $setup(posedge WDATA[9], posedge WCLKN, 1.0);
   $setup(negedge WDATA[9], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[9], 1.0);
   $hold(posedge WCLKN, negedge WDATA[9], 1.0);
   $setup(posedge WDATA[10], posedge WCLKN, 1.0);
   $setup(negedge WDATA[10], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[10], 1.0);
   $hold(posedge WCLKN, negedge WDATA[10], 1.0);
   $setup(posedge WDATA[11], posedge WCLKN, 1.0);
   $setup(negedge WDATA[11], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[11], 1.0);
   $hold(posedge WCLKN, negedge WDATA[11], 1.0);
   $setup(posedge WDATA[12], posedge WCLKN, 1.0);
   $setup(negedge WDATA[12], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[12], 1.0);
   $hold(posedge WCLKN, negedge WDATA[12], 1.0);
   $setup(posedge WDATA[13], posedge WCLKN, 1.0);
   $setup(negedge WDATA[13], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[13], 1.0);
   $hold(posedge WCLKN, negedge WDATA[13], 1.0);
   $setup(posedge WDATA[14], posedge WCLKN, 1.0);
   $setup(negedge WDATA[14], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[14], 1.0);
   $hold(posedge WCLKN, negedge WDATA[14], 1.0);
   $setup(posedge WDATA[15], posedge WCLKN, 1.0);
   $setup(negedge WDATA[15], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[15], 1.0);
   $hold(posedge WCLKN, negedge WDATA[15], 1.0);
   $setup(posedge WCLKE, posedge WCLKN, 1.0);
   $setup(negedge WCLKE, posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WCLKE, 1.0);
   $hold(posedge WCLKN, negedge WCLKE, 1.0);
   $setup(posedge WE, posedge WCLKN, 1.0);
   $setup(negedge WE, posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WE, 1.0);
   $hold(posedge WCLKN, negedge WE, 1.0);
   $setup(posedge RADDR[0], posedge RCLKN, 1.0);
   $setup(negedge RADDR[0], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[0], 1.0);
   $hold(posedge RCLKN, negedge RADDR[0], 1.0);
   $setup(posedge RADDR[1], posedge RCLKN, 1.0);
   $setup(negedge RADDR[1], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[1], 1.0);
   $hold(posedge RCLKN, negedge RADDR[1], 1.0);
   $setup(posedge RADDR[2], posedge RCLKN, 1.0);
   $setup(negedge RADDR[2], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[2], 1.0);
   $hold(posedge RCLKN, negedge RADDR[2], 1.0);
   $setup(posedge RADDR[3], posedge RCLKN, 1.0);
   $setup(negedge RADDR[3], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[3], 1.0);
   $hold(posedge RCLKN, negedge RADDR[3], 1.0);
   $setup(posedge RADDR[4], posedge RCLKN, 1.0);
   $setup(negedge RADDR[4], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[4], 1.0);
   $hold(posedge RCLKN, negedge RADDR[4], 1.0);
   $setup(posedge RADDR[5], posedge RCLKN, 1.0);
   $setup(negedge RADDR[5], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[5], 1.0);
   $hold(posedge RCLKN, negedge RADDR[5], 1.0);
   $setup(posedge RADDR[6], posedge RCLKN, 1.0);
   $setup(negedge RADDR[6], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[6], 1.0);
   $hold(posedge RCLKN, negedge RADDR[6], 1.0);
   $setup(posedge RADDR[7], posedge RCLKN, 1.0);
   $setup(negedge RADDR[7], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[7], 1.0);
   $hold(posedge RCLKN, negedge RADDR[7], 1.0);
   $setup(posedge RCLKE, posedge RCLKN, 1.0);
   $setup(negedge RCLKE, posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RCLKE, 1.0);
   $hold(posedge RCLKN, negedge RCLKE, 1.0);
   $setup(posedge RE, posedge RCLKN, 1.0);
   $setup(negedge RE, posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RE, 1.0);
   $hold(posedge RCLKN, negedge RE, 1.0);
   $recovery(posedge RCLKN, posedge WCLKN, 1.0);
   $recovery(negedge RCLKN, posedge WCLKN, 1.0);
   $removal(posedge RCLKN, posedge WCLKN, 1.0);
   $removal(negedge RCLKN, posedge WCLKN, 1.0);
   $recovery(posedge WCLKN, posedge RCLKN, 1.0);
   $recovery(negedge WCLKN, posedge RCLKN, 1.0);
   $removal(posedge WCLKN, posedge RCLKN, 1.0);
   $removal(negedge WCLKN, posedge RCLKN, 1.0);

endspecify
`endif

endmodule //SB_RAM4KNRNW



`timescale 1ps/1ps
module SB_RAM4K (RDATA, RCLK, RCLKE, RE, RADDR, WCLK, WCLKE, WE, WADDR, MASK, WDATA);
output [15:0] RDATA;
input RCLK;
input RCLKE;
input RE;
input [7:0] RADDR;
input WCLK;
input WCLKE;
input WE;
input [7:0] WADDR;
input [15:0] MASK;
input [15:0] WDATA;

assign (weak0, weak1) MASK = 16'b0;

parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

// local Parameters
localparam			CLOCK_PERIOD = 200;	//
localparam 			DELAY	= (CLOCK_PERIOD/10);		// Clock-to-output delay. Zero
							// time delays can be confusing
							// and sometimes cause problems.
localparam 			BUS_WIDTH = 16;		// Width of RAM (number of bits)

localparam 			ADDRESS_BUS_SIZE = 8;	// Number of bits required to
							// represent the RAM address

localparam   ADDRESSABLE_SPACE  = 2**ADDRESS_BUS_SIZE;	// Decimal address range [2^Size:0]


// SIGNAL DECLARATIONS
wire			   	WCLK_g, RCLK_g;
reg 				WCLKE_sync, RCLKE_sync; 
assign (weak0, weak1) RCLKE =1'b1 ;
assign (weak0, weak1) RE =1'b0 ;
assign (weak0, weak1) WCLKE =1'b1 ;
assign (weak0, weak1) WE =1'b0 ;
//reg  [BUS_WIDTH-1:0] Memory [ADDRESSABLE_SPACE-1:0];	// The RAM
reg	Memory	[BUS_WIDTH*ADDRESSABLE_SPACE-1:0];
// 
event Read_e, Write_e;

//////////////////// Collision detect begins here ///////////////////////////////
localparam 	TRUE = 1'b1;
localparam	FALSE = 1'b0;
reg 		Time_Collision_Detected = 1'b0;
wire		Address_Collision_Detected;

event Collision_e;

time COLLISION_TIME_WINDOW = (CLOCK_PERIOD/8); // This is an arbitray value, but is better than using an absolute 
						    // value, because the actual time window depends on the actual silicon 
						    // implementation. Thus the test is indicative of an Error and not
						    // guaranteed to be an error. Even so this is usefull.
time time_WCLK_RCLK, time_WCLK, time_RCLK;


//function reg Check_Timed_Window_Violation;
function	Check_Timed_Window_Violation;	//	by Jeffrey
input T1, T2, Minimum_Time_Window;
time T1, T2;
time Minimum_Time_Window;
time Difference;	
	begin
		Difference = (T1 - T2);
		if (Difference < 0) Difference = -Difference;
		Check_Timed_Window_Violation = (Difference < Minimum_Time_Window);
	end
endfunction


initial begin
       time_WCLK = CLOCK_PERIOD;	// Arbitrary initialisation value, ensure no window collison error on first clock edge.
       time_RCLK = (CLOCK_PERIOD*8);	// Arbitrary initialisation difference value, ensure no collision error on first clock edge.					
end

integer	i,j;

genvar k;
wire [7:0] RADDR_g;
wire [7:0] WADDR_g;
wire [15:0] WDATA_g;
for (k = 0; k < 8; k = k + 1) begin
	assign RADDR_g[k] = (RADDR[k] === 1'bz)? 1'b0 : RADDR[k];
	assign WADDR_g[k] = (WADDR[k] === 1'bz)? 1'b0 : WADDR[k];
	assign WDATA_g[k] = (WDATA[k] === 1'bz)? 1'b0 : WDATA[k];
	assign WDATA_g[k+8] = (WDATA[k+8] === 1'bz)? 1'b0 : WDATA[k+8];
end

initial	//	initialize ram_4k by parameter, section by section
begin
	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[BUS_WIDTH*i+j]	=	INIT_0[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*1+BUS_WIDTH*i+j]	=	INIT_1[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*2+BUS_WIDTH*i+j]	=	INIT_2[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*3+BUS_WIDTH*i+j]	=	INIT_3[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*4+BUS_WIDTH*i+j]	=	INIT_4[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*5+BUS_WIDTH*i+j]	=	INIT_5[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*6+BUS_WIDTH*i+j]	=	INIT_6[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*7+BUS_WIDTH*i+j]	=	INIT_7[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*8+BUS_WIDTH*i+j]	=	INIT_8[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*9+BUS_WIDTH*i+j]	=	INIT_9[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*10+BUS_WIDTH*i+j]	=	INIT_A[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*11+BUS_WIDTH*i+j]	=	INIT_B[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*12+BUS_WIDTH*i+j]	=	INIT_C[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*13+BUS_WIDTH*i+j]	=	INIT_D[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*14+BUS_WIDTH*i+j]	=	INIT_E[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*15+BUS_WIDTH*i+j]	=	INIT_F[BUS_WIDTH*i+j];
	end

end

assign Address_Collision_Detected = ((RE & WE & WCLKE & RCLKE)&(WADDR == RADDR)); 

always @(WCLK or WCLKE) 
begin 
	if(~WCLK)
	WCLKE_sync = WCLKE;   	
end 

always @(RCLK or RCLKE) 
begin 
	if (~RCLK)
	RCLKE_sync = RCLKE; 	
end 

assign WCLK_g = WCLK & WCLKE_sync;
assign RCLK_g = RCLK & RCLKE_sync;

always @(posedge WCLK_g) begin
	time_WCLK = $time;
end

always @(posedge RCLK_g) begin
    	time_RCLK = $time;
end
integer	SB_RAM4K_RDATA_log_file;									//.....................
initial	SB_RAM4K_RDATA_log_file=("SB_RAM4K_RDATA_log_file.txt");	//.....................
always @(posedge WCLK_g) begin

	Time_Collision_Detected = Check_Timed_Window_Violation(time_WCLK,time_RCLK,COLLISION_TIME_WINDOW);
        if (Time_Collision_Detected & Address_Collision_Detected)begin
        	$display("Warning: Write-Read collision detected, Data read value is XXXX\n");
 		$display("WCLK Time: %.3f   RCLK Time:%.3f  ",time_WCLK, time_RCLK,"WADDR: %d   RADDR:%d\n",WADDR, RADDR); 
 		$fdisplay(SB_RAM4K_RDATA_log_file,"Warning: Write-Read collision detected, Data read value is XXXX\n");
		$fdisplay(SB_RAM4K_RDATA_log_file,"WCLK Time: %.3f   RCLK Time:%.3f  ",time_WCLK, time_RCLK, "WADDR: %d   RADDR:%d\n",WADDR, RADDR); 	
 		-> Collision_e;
	end
end




//	code modify for universal verilog compiler

always @ (posedge WCLK_g)
begin
	if	(WE)
	begin
		-> Write_e;
		for	(i=0;i<=BUS_WIDTH-1; i=i+1)
		begin
			if	(MASK[i] !=1)
				Memory[WADDR_g*BUS_WIDTH+i]	<=	WDATA_g[i];
			else
				Memory[WADDR_g*BUS_WIDTH+i]	<=	Memory[WADDR_g*BUS_WIDTH+i];
		end
	end
end

//reg	[15:0]	RDATA = 0;
reg	[15:0]	RDATA;

initial
begin
   RDATA = $random;
end

// Look at the rising edge of the clock

always @ (posedge RCLK_g)
begin
	if	(RE)
	begin
		-> Read_e;
		if	(Time_Collision_Detected & Address_Collision_Detected) 
			RDATA <= 16'hXXXX;
		else
			for	(i=0;i<=BUS_WIDTH-1;i=i+1)
				RDATA[i]	<= Memory[RADDR_g*BUS_WIDTH+i];
	end
end

`ifdef TIMINGCHECK
specify
   (RCLK *> RDATA[0]) = (1.0, 1.0);
   (RCLK *> RDATA[1]) = (1.0, 1.0);
   (RCLK *> RDATA[2]) = (1.0, 1.0);
   (RCLK *> RDATA[3]) = (1.0, 1.0);
   (RCLK *> RDATA[4]) = (1.0, 1.0);
   (RCLK *> RDATA[5]) = (1.0, 1.0);
   (RCLK *> RDATA[6]) = (1.0, 1.0);
   (RCLK *> RDATA[7]) = (1.0, 1.0);
   (RCLK *> RDATA[8]) = (1.0, 1.0);
   (RCLK *> RDATA[9]) = (1.0, 1.0);
   (RCLK *> RDATA[10]) = (1.0, 1.0);
   (RCLK *> RDATA[11]) = (1.0, 1.0);
   (RCLK *> RDATA[12]) = (1.0, 1.0);
   (RCLK *> RDATA[13]) = (1.0, 1.0);
   (RCLK *> RDATA[14]) = (1.0, 1.0);
   (RCLK *> RDATA[15]) = (1.0, 1.0);
   $setup(posedge MASK[0], posedge WCLK, 1.0);
   $setup(negedge MASK[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[0], 1.0);
   $hold(posedge WCLK, negedge MASK[0], 1.0);
   $setup(posedge MASK[1], posedge WCLK, 1.0);
   $setup(negedge MASK[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[1], 1.0);
   $hold(posedge WCLK, negedge MASK[1], 1.0);
   $setup(posedge MASK[2], posedge WCLK, 1.0);
   $setup(negedge MASK[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[2], 1.0);
   $hold(posedge WCLK, negedge MASK[2], 1.0);
   $setup(posedge MASK[3], posedge WCLK, 1.0);
   $setup(negedge MASK[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[3], 1.0);
   $hold(posedge WCLK, negedge MASK[3], 1.0);
   $setup(posedge MASK[4], posedge WCLK, 1.0);
   $setup(negedge MASK[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[4], 1.0);
   $hold(posedge WCLK, negedge MASK[4], 1.0);
   $setup(posedge MASK[5], posedge WCLK, 1.0);
   $setup(negedge MASK[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[5], 1.0);
   $hold(posedge WCLK, negedge MASK[5], 1.0);
   $setup(posedge MASK[6], posedge WCLK, 1.0);
   $setup(negedge MASK[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[6], 1.0);
   $hold(posedge WCLK, negedge MASK[6], 1.0);
   $setup(posedge MASK[7], posedge WCLK, 1.0);
   $setup(negedge MASK[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[7], 1.0);
   $hold(posedge WCLK, negedge MASK[7], 1.0);
   $setup(posedge MASK[8], posedge WCLK, 1.0);
   $setup(negedge MASK[8], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[8], 1.0);
   $hold(posedge WCLK, negedge MASK[8], 1.0);
   $setup(posedge MASK[9], posedge WCLK, 1.0);
   $setup(negedge MASK[9], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[9], 1.0);
   $hold(posedge WCLK, negedge MASK[9], 1.0);
   $setup(posedge MASK[10], posedge WCLK, 1.0);
   $setup(negedge MASK[10], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[10], 1.0);
   $hold(posedge WCLK, negedge MASK[10], 1.0);
   $setup(posedge MASK[11], posedge WCLK, 1.0);
   $setup(negedge MASK[11], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[11], 1.0);
   $hold(posedge WCLK, negedge MASK[11], 1.0);
   $setup(posedge MASK[12], posedge WCLK, 1.0);
   $setup(negedge MASK[12], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[12], 1.0);
   $hold(posedge WCLK, negedge MASK[12], 1.0);
   $setup(posedge MASK[13], posedge WCLK, 1.0);
   $setup(negedge MASK[13], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[13], 1.0);
   $hold(posedge WCLK, negedge MASK[13], 1.0);
   $setup(posedge MASK[14], posedge WCLK, 1.0);
   $setup(negedge MASK[14], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[14], 1.0);
   $hold(posedge WCLK, negedge MASK[14], 1.0);
   $setup(posedge MASK[15], posedge WCLK, 1.0);
   $setup(negedge MASK[15], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[15], 1.0);
   $hold(posedge WCLK, negedge MASK[15], 1.0);
   $setup(posedge WADDR[0], posedge WCLK, 1.0);
   $setup(negedge WADDR[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[0], 1.0);
   $hold(posedge WCLK, negedge WADDR[0], 1.0);
   $setup(posedge WADDR[1], posedge WCLK, 1.0);
   $setup(negedge WADDR[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[1], 1.0);
   $hold(posedge WCLK, negedge WADDR[1], 1.0);
   $setup(posedge WADDR[2], posedge WCLK, 1.0);
   $setup(negedge WADDR[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[2], 1.0);
   $hold(posedge WCLK, negedge WADDR[2], 1.0);
   $setup(posedge WADDR[3], posedge WCLK, 1.0);
   $setup(negedge WADDR[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[3], 1.0);
   $hold(posedge WCLK, negedge WADDR[3], 1.0);
   $setup(posedge WADDR[4], posedge WCLK, 1.0);
   $setup(negedge WADDR[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[4], 1.0);
   $hold(posedge WCLK, negedge WADDR[4], 1.0);
   $setup(posedge WADDR[5], posedge WCLK, 1.0);
   $setup(negedge WADDR[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[5], 1.0);
   $hold(posedge WCLK, negedge WADDR[5], 1.0);
   $setup(posedge WADDR[6], posedge WCLK, 1.0);
   $setup(negedge WADDR[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[6], 1.0);
   $hold(posedge WCLK, negedge WADDR[6], 1.0);
   $setup(posedge WADDR[7], posedge WCLK, 1.0);
   $setup(negedge WADDR[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[7], 1.0);
   $hold(posedge WCLK, negedge WADDR[7], 1.0);
   $setup(posedge WDATA[0], posedge WCLK, 1.0);
   $setup(negedge WDATA[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[0], 1.0);
   $hold(posedge WCLK, negedge WDATA[0], 1.0);
   $setup(posedge WDATA[1], posedge WCLK, 1.0);
   $setup(negedge WDATA[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[1], 1.0);
   $hold(posedge WCLK, negedge WDATA[1], 1.0);
   $setup(posedge WDATA[2], posedge WCLK, 1.0);
   $setup(negedge WDATA[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[2], 1.0);
   $hold(posedge WCLK, negedge WDATA[2], 1.0);
   $setup(posedge WDATA[3], posedge WCLK, 1.0);
   $setup(negedge WDATA[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[3], 1.0);
   $hold(posedge WCLK, negedge WDATA[3], 1.0);
   $setup(posedge WDATA[4], posedge WCLK, 1.0);
   $setup(negedge WDATA[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[4], 1.0);
   $hold(posedge WCLK, negedge WDATA[4], 1.0);
   $setup(posedge WDATA[5], posedge WCLK, 1.0);
   $setup(negedge WDATA[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[5], 1.0);
   $hold(posedge WCLK, negedge WDATA[5], 1.0);
   $setup(posedge WDATA[6], posedge WCLK, 1.0);
   $setup(negedge WDATA[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[6], 1.0);
   $hold(posedge WCLK, negedge WDATA[6], 1.0);
   $setup(posedge WDATA[7], posedge WCLK, 1.0);
   $setup(negedge WDATA[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[7], 1.0);
   $hold(posedge WCLK, negedge WDATA[7], 1.0);
   $setup(posedge WDATA[8], posedge WCLK, 1.0);
   $setup(negedge WDATA[8], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[8], 1.0);
   $hold(posedge WCLK, negedge WDATA[8], 1.0);
   $setup(posedge WDATA[9], posedge WCLK, 1.0);
   $setup(negedge WDATA[9], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[9], 1.0);
   $hold(posedge WCLK, negedge WDATA[9], 1.0);
   $setup(posedge WDATA[10], posedge WCLK, 1.0);
   $setup(negedge WDATA[10], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[10], 1.0);
   $hold(posedge WCLK, negedge WDATA[10], 1.0);
   $setup(posedge WDATA[11], posedge WCLK, 1.0);
   $setup(negedge WDATA[11], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[11], 1.0);
   $hold(posedge WCLK, negedge WDATA[11], 1.0);
   $setup(posedge WDATA[12], posedge WCLK, 1.0);
   $setup(negedge WDATA[12], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[12], 1.0);
   $hold(posedge WCLK, negedge WDATA[12], 1.0);
   $setup(posedge WDATA[13], posedge WCLK, 1.0);
   $setup(negedge WDATA[13], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[13], 1.0);
   $hold(posedge WCLK, negedge WDATA[13], 1.0);
   $setup(posedge WDATA[14], posedge WCLK, 1.0);
   $setup(negedge WDATA[14], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[14], 1.0);
   $hold(posedge WCLK, negedge WDATA[14], 1.0);
   $setup(posedge WDATA[15], posedge WCLK, 1.0);
   $setup(negedge WDATA[15], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[15], 1.0);
   $hold(posedge WCLK, negedge WDATA[15], 1.0);
   $setup(posedge WCLKE, posedge WCLK, 1.0);
   $setup(negedge WCLKE, posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WCLKE, 1.0);
   $hold(posedge WCLK, negedge WCLKE, 1.0);
   $setup(posedge WE, posedge WCLK, 1.0);
   $setup(negedge WE, posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WE, 1.0);
   $hold(posedge WCLK, negedge WE, 1.0);
   $setup(posedge RADDR[0], posedge RCLK, 1.0);
   $setup(negedge RADDR[0], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[0], 1.0);
   $hold(posedge RCLK, negedge RADDR[0], 1.0);
   $setup(posedge RADDR[1], posedge RCLK, 1.0);
   $setup(negedge RADDR[1], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[1], 1.0);
   $hold(posedge RCLK, negedge RADDR[1], 1.0);
   $setup(posedge RADDR[2], posedge RCLK, 1.0);
   $setup(negedge RADDR[2], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[2], 1.0);
   $hold(posedge RCLK, negedge RADDR[2], 1.0);
   $setup(posedge RADDR[3], posedge RCLK, 1.0);
   $setup(negedge RADDR[3], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[3], 1.0);
   $hold(posedge RCLK, negedge RADDR[3], 1.0);
   $setup(posedge RADDR[4], posedge RCLK, 1.0);
   $setup(negedge RADDR[4], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[4], 1.0);
   $hold(posedge RCLK, negedge RADDR[4], 1.0);
   $setup(posedge RADDR[5], posedge RCLK, 1.0);
   $setup(negedge RADDR[5], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[5], 1.0);
   $hold(posedge RCLK, negedge RADDR[5], 1.0);
   $setup(posedge RADDR[6], posedge RCLK, 1.0);
   $setup(negedge RADDR[6], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[6], 1.0);
   $hold(posedge RCLK, negedge RADDR[6], 1.0);
   $setup(posedge RADDR[7], posedge RCLK, 1.0);
   $setup(negedge RADDR[7], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[7], 1.0);
   $hold(posedge RCLK, negedge RADDR[7], 1.0);
   $setup(posedge RCLKE, posedge RCLK, 1.0);
   $setup(negedge RCLKE, posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RCLKE, 1.0);
   $hold(posedge RCLK, negedge RCLKE, 1.0);
   $setup(posedge RE, posedge RCLK, 1.0);
   $setup(negedge RE, posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RE, 1.0);
   $hold(posedge RCLK, negedge RE, 1.0);
   // $recovery(posedge RCLK, posedge WCLK, 1.0);
   // $recovery(negedge RCLK, posedge WCLK, 1.0);
   // $removal(posedge RCLK, posedge WCLK, 1.0);
   // $removal(negedge RCLK, posedge WCLK, 1.0);
   // $recovery(posedge WCLK, posedge RCLK, 1.0);
   // $recovery(negedge WCLK, posedge RCLK, 1.0);
   // $removal(posedge WCLK, posedge RCLK, 1.0);
   // $removal(negedge WCLK, posedge RCLK, 1.0);

endspecify
`endif

endmodule	 //	SB_RAM4K


/*****ice40P08 RAM prims******/
`timescale 1ps/1ps
module SB_RAM40_4KNR (RDATA, RCLKN, RCLKE, RE, RADDR, WCLK, WCLKE, WE, WADDR, MASK, WDATA);
output [15:0] RDATA;
input RCLKN;
input RCLKE;
input RE;
input [10:0] RADDR;
input WCLK;
input WCLKE;
input WE;
input [10:0] WADDR;
input [15:0] MASK;
input [15:0] WDATA;

parameter WRITE_MODE = 0; /// can be integer 0(256X16 mode) or 1(512X8 mode) or 2(1024X4 mode) or 3(2048X2 mode)
parameter READ_MODE = 0;  /// can be integer 0(256X16 mode) or 1(512X8 mode) or 2(1024X4 mode) or 3(2048X2 mode)


parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

wire RCLK;
assign (weak0, weak1) RCLKE =1'b1 ;
assign (weak0, weak1) RE =1'b0 ;
assign (weak0, weak1) WCLKE =1'b1 ;
assign (weak0, weak1) WE =1'b0 ;
assign RCLK = ~RCLKN;

SB_RAM40_4K ram40_4K_nr_inst (
	.RDATA(RDATA),
	.RCLK(RCLK),
	.RCLKE(RCLKE),
	.RE(RE),
	.RADDR(RADDR),
	.WCLK(WCLK),
	.WCLKE(WCLKE),
	.WE(WE),
	.WADDR(WADDR),
	.MASK(MASK),
	.WDATA(WDATA));

defparam ram40_4K_nr_inst.WRITE_MODE = WRITE_MODE;
defparam ram40_4K_nr_inst.READ_MODE = READ_MODE;
defparam ram40_4K_nr_inst.INIT_0 = INIT_0;
defparam ram40_4K_nr_inst.INIT_1 = INIT_1;
defparam ram40_4K_nr_inst.INIT_2 = INIT_2;
defparam ram40_4K_nr_inst.INIT_3 = INIT_3;
defparam ram40_4K_nr_inst.INIT_4 = INIT_4;
defparam ram40_4K_nr_inst.INIT_5 = INIT_5;
defparam ram40_4K_nr_inst.INIT_6 = INIT_6;
defparam ram40_4K_nr_inst.INIT_7 = INIT_7;
defparam ram40_4K_nr_inst.INIT_8 = INIT_8;
defparam ram40_4K_nr_inst.INIT_9 = INIT_9;
defparam ram40_4K_nr_inst.INIT_A = INIT_A;
defparam ram40_4K_nr_inst.INIT_B = INIT_B;
defparam ram40_4K_nr_inst.INIT_C = INIT_C;
defparam ram40_4K_nr_inst.INIT_D = INIT_D;
defparam ram40_4K_nr_inst.INIT_E = INIT_E;
defparam ram40_4K_nr_inst.INIT_F = INIT_F;

`ifdef TIMINGCHECK
specify
   (RCLKN *> RDATA[0]) = (1.0, 1.0);
   (RCLKN *> RDATA[1]) = (1.0, 1.0);
   (RCLKN *> RDATA[2]) = (1.0, 1.0);
   (RCLKN *> RDATA[3]) = (1.0, 1.0);
   (RCLKN *> RDATA[4]) = (1.0, 1.0);
   (RCLKN *> RDATA[5]) = (1.0, 1.0);
   (RCLKN *> RDATA[6]) = (1.0, 1.0);
   (RCLKN *> RDATA[7]) = (1.0, 1.0);
   (RCLKN *> RDATA[8]) = (1.0, 1.0);
   (RCLKN *> RDATA[9]) = (1.0, 1.0);
   (RCLKN *> RDATA[10]) = (1.0, 1.0);
   (RCLKN *> RDATA[11]) = (1.0, 1.0);
   (RCLKN *> RDATA[12]) = (1.0, 1.0);
   (RCLKN *> RDATA[13]) = (1.0, 1.0);
   (RCLKN *> RDATA[14]) = (1.0, 1.0);
   (RCLKN *> RDATA[15]) = (1.0, 1.0);
   $setup(posedge MASK[0], posedge WCLK, 1.0);
   $setup(negedge MASK[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[0], 1.0);
   $hold(posedge WCLK, negedge MASK[0], 1.0);
   $setup(posedge MASK[1], posedge WCLK, 1.0);
   $setup(negedge MASK[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[1], 1.0);
   $hold(posedge WCLK, negedge MASK[1], 1.0);
   $setup(posedge MASK[2], posedge WCLK, 1.0);
   $setup(negedge MASK[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[2], 1.0);
   $hold(posedge WCLK, negedge MASK[2], 1.0);
   $setup(posedge MASK[3], posedge WCLK, 1.0);
   $setup(negedge MASK[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[3], 1.0);
   $hold(posedge WCLK, negedge MASK[3], 1.0);
   $setup(posedge MASK[4], posedge WCLK, 1.0);
   $setup(negedge MASK[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[4], 1.0);
   $hold(posedge WCLK, negedge MASK[4], 1.0);
   $setup(posedge MASK[5], posedge WCLK, 1.0);
   $setup(negedge MASK[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[5], 1.0);
   $hold(posedge WCLK, negedge MASK[5], 1.0);
   $setup(posedge MASK[6], posedge WCLK, 1.0);
   $setup(negedge MASK[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[6], 1.0);
   $hold(posedge WCLK, negedge MASK[6], 1.0);
   $setup(posedge MASK[7], posedge WCLK, 1.0);
   $setup(negedge MASK[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[7], 1.0);
   $hold(posedge WCLK, negedge MASK[7], 1.0);
   $setup(posedge MASK[8], posedge WCLK, 1.0);
   $setup(negedge MASK[8], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[8], 1.0);
   $hold(posedge WCLK, negedge MASK[8], 1.0);
   $setup(posedge MASK[9], posedge WCLK, 1.0);
   $setup(negedge MASK[9], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[9], 1.0);
   $hold(posedge WCLK, negedge MASK[9], 1.0);
   $setup(posedge MASK[10], posedge WCLK, 1.0);
   $setup(negedge MASK[10], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[10], 1.0);
   $hold(posedge WCLK, negedge MASK[10], 1.0);
   $setup(posedge MASK[11], posedge WCLK, 1.0);
   $setup(negedge MASK[11], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[11], 1.0);
   $hold(posedge WCLK, negedge MASK[11], 1.0);
   $setup(posedge MASK[12], posedge WCLK, 1.0);
   $setup(negedge MASK[12], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[12], 1.0);
   $hold(posedge WCLK, negedge MASK[12], 1.0);
   $setup(posedge MASK[13], posedge WCLK, 1.0);
   $setup(negedge MASK[13], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[13], 1.0);
   $hold(posedge WCLK, negedge MASK[13], 1.0);
   $setup(posedge MASK[14], posedge WCLK, 1.0);
   $setup(negedge MASK[14], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[14], 1.0);
   $hold(posedge WCLK, negedge MASK[14], 1.0);
   $setup(posedge MASK[15], posedge WCLK, 1.0);
   $setup(negedge MASK[15], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[15], 1.0);
   $hold(posedge WCLK, negedge MASK[15], 1.0);
   $setup(posedge WADDR[0], posedge WCLK, 1.0);
   $setup(negedge WADDR[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[0], 1.0);
   $hold(posedge WCLK, negedge WADDR[0], 1.0);
   $setup(posedge WADDR[1], posedge WCLK, 1.0);
   $setup(negedge WADDR[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[1], 1.0);
   $hold(posedge WCLK, negedge WADDR[1], 1.0);
   $setup(posedge WADDR[2], posedge WCLK, 1.0);
   $setup(negedge WADDR[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[2], 1.0);
   $hold(posedge WCLK, negedge WADDR[2], 1.0);
   $setup(posedge WADDR[3], posedge WCLK, 1.0);
   $setup(negedge WADDR[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[3], 1.0);
   $hold(posedge WCLK, negedge WADDR[3], 1.0);
   $setup(posedge WADDR[4], posedge WCLK, 1.0);
   $setup(negedge WADDR[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[4], 1.0);
   $hold(posedge WCLK, negedge WADDR[4], 1.0);
   $setup(posedge WADDR[5], posedge WCLK, 1.0);
   $setup(negedge WADDR[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[5], 1.0);
   $hold(posedge WCLK, negedge WADDR[5], 1.0);
   $setup(posedge WADDR[6], posedge WCLK, 1.0);
   $setup(negedge WADDR[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[6], 1.0);
   $hold(posedge WCLK, negedge WADDR[6], 1.0);
   $setup(posedge WADDR[7], posedge WCLK, 1.0);
   $setup(negedge WADDR[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[7], 1.0);
   $hold(posedge WCLK, negedge WADDR[7], 1.0);
   $setup(posedge WADDR[8], posedge WCLK, 1.0);
   $setup(negedge WADDR[8], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[8], 1.0);
   $hold(posedge WCLK, negedge WADDR[8], 1.0);
   $setup(posedge WADDR[9], posedge WCLK, 1.0);
   $setup(negedge WADDR[9], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[9], 1.0);
   $hold(posedge WCLK, negedge WADDR[9], 1.0);
   $setup(posedge WADDR[10], posedge WCLK, 1.0);
   $setup(negedge WADDR[10], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[10], 1.0);
   $hold(posedge WCLK, negedge WADDR[10], 1.0);
   $setup(posedge WDATA[0], posedge WCLK, 1.0);
   $setup(negedge WDATA[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[0], 1.0);
   $hold(posedge WCLK, negedge WDATA[0], 1.0);
   $setup(posedge WDATA[1], posedge WCLK, 1.0);
   $setup(negedge WDATA[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[1], 1.0);
   $hold(posedge WCLK, negedge WDATA[1], 1.0);
   $setup(posedge WDATA[2], posedge WCLK, 1.0);
   $setup(negedge WDATA[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[2], 1.0);
   $hold(posedge WCLK, negedge WDATA[2], 1.0);
   $setup(posedge WDATA[3], posedge WCLK, 1.0);
   $setup(negedge WDATA[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[3], 1.0);
   $hold(posedge WCLK, negedge WDATA[3], 1.0);
   $setup(posedge WDATA[4], posedge WCLK, 1.0);
   $setup(negedge WDATA[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[4], 1.0);
   $hold(posedge WCLK, negedge WDATA[4], 1.0);
   $setup(posedge WDATA[5], posedge WCLK, 1.0);
   $setup(negedge WDATA[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[5], 1.0);
   $hold(posedge WCLK, negedge WDATA[5], 1.0);
   $setup(posedge WDATA[6], posedge WCLK, 1.0);
   $setup(negedge WDATA[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[6], 1.0);
   $hold(posedge WCLK, negedge WDATA[6], 1.0);
   $setup(posedge WDATA[7], posedge WCLK, 1.0);
   $setup(negedge WDATA[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[7], 1.0);
   $hold(posedge WCLK, negedge WDATA[7], 1.0);
   $setup(posedge WDATA[8], posedge WCLK, 1.0);
   $setup(negedge WDATA[8], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[8], 1.0);
   $hold(posedge WCLK, negedge WDATA[8], 1.0);
   $setup(posedge WDATA[9], posedge WCLK, 1.0);
   $setup(negedge WDATA[9], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[9], 1.0);
   $hold(posedge WCLK, negedge WDATA[9], 1.0);
   $setup(posedge WDATA[10], posedge WCLK, 1.0);
   $setup(negedge WDATA[10], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[10], 1.0);
   $hold(posedge WCLK, negedge WDATA[10], 1.0);
   $setup(posedge WDATA[11], posedge WCLK, 1.0);
   $setup(negedge WDATA[11], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[11], 1.0);
   $hold(posedge WCLK, negedge WDATA[11], 1.0);
   $setup(posedge WDATA[12], posedge WCLK, 1.0);
   $setup(negedge WDATA[12], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[12], 1.0);
   $hold(posedge WCLK, negedge WDATA[12], 1.0);
   $setup(posedge WDATA[13], posedge WCLK, 1.0);
   $setup(negedge WDATA[13], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[13], 1.0);
   $hold(posedge WCLK, negedge WDATA[13], 1.0);
   $setup(posedge WDATA[14], posedge WCLK, 1.0);
   $setup(negedge WDATA[14], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[14], 1.0);
   $hold(posedge WCLK, negedge WDATA[14], 1.0);
   $setup(posedge WDATA[15], posedge WCLK, 1.0);
   $setup(negedge WDATA[15], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[15], 1.0);
   $hold(posedge WCLK, negedge WDATA[15], 1.0);
   $setup(posedge WCLKE, posedge WCLK, 1.0);
   $setup(negedge WCLKE, posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WCLKE, 1.0);
   $hold(posedge WCLK, negedge WCLKE, 1.0);
   $setup(posedge WE, posedge WCLK, 1.0);
   $setup(negedge WE, posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WE, 1.0);
   $hold(posedge WCLK, negedge WE, 1.0);
   $setup(posedge RADDR[0], posedge RCLKN, 1.0);
   $setup(negedge RADDR[0], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[0], 1.0);
   $hold(posedge RCLKN, negedge RADDR[0], 1.0);
   $setup(posedge RADDR[1], posedge RCLKN, 1.0);
   $setup(negedge RADDR[1], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[1], 1.0);
   $hold(posedge RCLKN, negedge RADDR[1], 1.0);
   $setup(posedge RADDR[2], posedge RCLKN, 1.0);
   $setup(negedge RADDR[2], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[2], 1.0);
   $hold(posedge RCLKN, negedge RADDR[2], 1.0);
   $setup(posedge RADDR[3], posedge RCLKN, 1.0);
   $setup(negedge RADDR[3], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[3], 1.0);
   $hold(posedge RCLKN, negedge RADDR[3], 1.0);
   $setup(posedge RADDR[4], posedge RCLKN, 1.0);
   $setup(negedge RADDR[4], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[4], 1.0);
   $hold(posedge RCLKN, negedge RADDR[4], 1.0);
   $setup(posedge RADDR[5], posedge RCLKN, 1.0);
   $setup(negedge RADDR[5], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[5], 1.0);
   $hold(posedge RCLKN, negedge RADDR[5], 1.0);
   $setup(posedge RADDR[6], posedge RCLKN, 1.0);
   $setup(negedge RADDR[6], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[6], 1.0);
   $hold(posedge RCLKN, negedge RADDR[6], 1.0);
   $setup(posedge RADDR[7], posedge RCLKN, 1.0);
   $setup(negedge RADDR[7], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[7], 1.0);
   $hold(posedge RCLKN, negedge RADDR[7], 1.0);
   $setup(posedge RADDR[8], posedge RCLKN, 1.0);
   $setup(negedge RADDR[8], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[8], 1.0);
   $hold(posedge RCLKN, negedge RADDR[8], 1.0);
   $setup(posedge RADDR[9], posedge RCLKN, 1.0);
   $setup(negedge RADDR[9], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[9], 1.0);
   $hold(posedge RCLKN, negedge RADDR[9], 1.0);
   $setup(posedge RADDR[10], posedge RCLKN, 1.0);
   $setup(negedge RADDR[10], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[10], 1.0);
   $hold(posedge RCLKN, negedge RADDR[10], 1.0);
   $setup(posedge RCLKE, posedge RCLKN, 1.0);
   $setup(negedge RCLKE, posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RCLKE, 1.0);
   $hold(posedge RCLKN, negedge RCLKE, 1.0);
   $setup(posedge RE, posedge RCLKN, 1.0);
   $setup(negedge RE, posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RE, 1.0);
   $hold(posedge RCLKN, negedge RE, 1.0);

endspecify
`endif

endmodule //SB_RAM40_4KNR

`timescale 1ps/1ps
module SB_RAM40_4KNW (RDATA, RCLK, RCLKE, RE, RADDR, WCLKN, WCLKE, WE, WADDR, MASK, WDATA);
output [15:0] RDATA;
input RCLK;
input RCLKE;
input RE;
input [10:0] RADDR;
input WCLKN;
input WCLKE;
input WE;
input [10:0] WADDR;
input [15:0] MASK;
input [15:0] WDATA;

parameter WRITE_MODE = 0; /// can be integer 0(256X16 mode) or 1(512X8 mode) or 2(1024X4 mode) or 3(2048X2 mode)
parameter READ_MODE = 0;  /// can be integer 0(256X16 mode) or 1(512X8 mode) or 2(1024X4 mode) or 3(2048X2 mode)


parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

wire WCLK;
assign (weak0, weak1) RCLKE =1'b1 ;
assign (weak0, weak1) RE =1'b0 ;
assign (weak0, weak1) WCLKE =1'b1 ;
assign (weak0, weak1) WE =1'b0 ;
assign WCLK = ~WCLKN;

SB_RAM40_4K ram40_4K_nw_inst (
	.RDATA(RDATA),
	.RCLK(RCLK),
	.RCLKE(RCLKE),
	.RE(RE),
	.RADDR(RADDR),
	.WCLK(WCLK),
	.WCLKE(WCLKE),
	.WE(WE),
	.WADDR(WADDR),
	.MASK(MASK),
	.WDATA(WDATA));

defparam ram40_4K_nw_inst.WRITE_MODE = WRITE_MODE;
defparam ram40_4K_nw_inst.READ_MODE = READ_MODE;
defparam ram40_4K_nw_inst.INIT_0 = INIT_0;
defparam ram40_4K_nw_inst.INIT_1 = INIT_1;
defparam ram40_4K_nw_inst.INIT_2 = INIT_2;
defparam ram40_4K_nw_inst.INIT_3 = INIT_3;
defparam ram40_4K_nw_inst.INIT_4 = INIT_4;
defparam ram40_4K_nw_inst.INIT_5 = INIT_5;
defparam ram40_4K_nw_inst.INIT_6 = INIT_6;
defparam ram40_4K_nw_inst.INIT_7 = INIT_7;
defparam ram40_4K_nw_inst.INIT_8 = INIT_8;
defparam ram40_4K_nw_inst.INIT_9 = INIT_9;
defparam ram40_4K_nw_inst.INIT_A = INIT_A;
defparam ram40_4K_nw_inst.INIT_B = INIT_B;
defparam ram40_4K_nw_inst.INIT_C = INIT_C;
defparam ram40_4K_nw_inst.INIT_D = INIT_D;
defparam ram40_4K_nw_inst.INIT_E = INIT_E;
defparam ram40_4K_nw_inst.INIT_F = INIT_F;


`ifdef TIMINGCHECK
specify
   (RCLK *> RDATA[0]) = (1.0, 1.0);
   (RCLK *> RDATA[1]) = (1.0, 1.0);
   (RCLK *> RDATA[2]) = (1.0, 1.0);
   (RCLK *> RDATA[3]) = (1.0, 1.0);
   (RCLK *> RDATA[4]) = (1.0, 1.0);
   (RCLK *> RDATA[5]) = (1.0, 1.0);
   (RCLK *> RDATA[6]) = (1.0, 1.0);
   (RCLK *> RDATA[7]) = (1.0, 1.0);
   (RCLK *> RDATA[8]) = (1.0, 1.0);
   (RCLK *> RDATA[9]) = (1.0, 1.0);
   (RCLK *> RDATA[10]) = (1.0, 1.0);
   (RCLK *> RDATA[11]) = (1.0, 1.0);
   (RCLK *> RDATA[12]) = (1.0, 1.0);
   (RCLK *> RDATA[13]) = (1.0, 1.0);
   (RCLK *> RDATA[14]) = (1.0, 1.0);
   (RCLK *> RDATA[15]) = (1.0, 1.0);
   $setup(posedge MASK[0], posedge WCLKN, 1.0);
   $setup(negedge MASK[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[0], 1.0);
   $hold(posedge WCLKN, negedge MASK[0], 1.0);
   $setup(posedge MASK[1], posedge WCLKN, 1.0);
   $setup(negedge MASK[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[1], 1.0);
   $hold(posedge WCLKN, negedge MASK[1], 1.0);
   $setup(posedge MASK[2], posedge WCLKN, 1.0);
   $setup(negedge MASK[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[2], 1.0);
   $hold(posedge WCLKN, negedge MASK[2], 1.0);
   $setup(posedge MASK[3], posedge WCLKN, 1.0);
   $setup(negedge MASK[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[3], 1.0);
   $hold(posedge WCLKN, negedge MASK[3], 1.0);
   $setup(posedge MASK[4], posedge WCLKN, 1.0);
   $setup(negedge MASK[4], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[4], 1.0);
   $hold(posedge WCLKN, negedge MASK[4], 1.0);
   $setup(posedge MASK[5], posedge WCLKN, 1.0);
   $setup(negedge MASK[5], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[5], 1.0);
   $hold(posedge WCLKN, negedge MASK[5], 1.0);
   $setup(posedge MASK[6], posedge WCLKN, 1.0);
   $setup(negedge MASK[6], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[6], 1.0);
   $hold(posedge WCLKN, negedge MASK[6], 1.0);
   $setup(posedge MASK[7], posedge WCLKN, 1.0);
   $setup(negedge MASK[7], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[7], 1.0);
   $hold(posedge WCLKN, negedge MASK[7], 1.0);
   $setup(posedge MASK[8], posedge WCLKN, 1.0);
   $setup(negedge MASK[8], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[8], 1.0);
   $hold(posedge WCLKN, negedge MASK[8], 1.0);
   $setup(posedge MASK[9], posedge WCLKN, 1.0);
   $setup(negedge MASK[9], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[9], 1.0);
   $hold(posedge WCLKN, negedge MASK[9], 1.0);
   $setup(posedge MASK[10], posedge WCLKN, 1.0);
   $setup(negedge MASK[10], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[10], 1.0);
   $hold(posedge WCLKN, negedge MASK[10], 1.0);
   $setup(posedge MASK[11], posedge WCLKN, 1.0);
   $setup(negedge MASK[11], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[11], 1.0);
   $hold(posedge WCLKN, negedge MASK[11], 1.0);
   $setup(posedge MASK[12], posedge WCLKN, 1.0);
   $setup(negedge MASK[12], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[12], 1.0);
   $hold(posedge WCLKN, negedge MASK[12], 1.0);
   $setup(posedge MASK[13], posedge WCLKN, 1.0);
   $setup(negedge MASK[13], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[13], 1.0);
   $hold(posedge WCLKN, negedge MASK[13], 1.0);
   $setup(posedge MASK[14], posedge WCLKN, 1.0);
   $setup(negedge MASK[14], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[14], 1.0);
   $hold(posedge WCLKN, negedge MASK[14], 1.0);
   $setup(posedge MASK[15], posedge WCLKN, 1.0);
   $setup(negedge MASK[15], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[15], 1.0);
   $hold(posedge WCLKN, negedge MASK[15], 1.0);
   $setup(posedge WADDR[0], posedge WCLKN, 1.0);
   $setup(negedge WADDR[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[0], 1.0);
   $hold(posedge WCLKN, negedge WADDR[0], 1.0);
   $setup(posedge WADDR[1], posedge WCLKN, 1.0);
   $setup(negedge WADDR[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[1], 1.0);
   $hold(posedge WCLKN, negedge WADDR[1], 1.0);
   $setup(posedge WADDR[2], posedge WCLKN, 1.0);
   $setup(negedge WADDR[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[2], 1.0);
   $hold(posedge WCLKN, negedge WADDR[2], 1.0);
   $setup(posedge WADDR[3], posedge WCLKN, 1.0);
   $setup(negedge WADDR[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[3], 1.0);
   $hold(posedge WCLKN, negedge WADDR[3], 1.0);
   $setup(posedge WADDR[4], posedge WCLKN, 1.0);
   $setup(negedge WADDR[4], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[4], 1.0);
   $hold(posedge WCLKN, negedge WADDR[4], 1.0);
   $setup(posedge WADDR[5], posedge WCLKN, 1.0);
   $setup(negedge WADDR[5], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[5], 1.0);
   $hold(posedge WCLKN, negedge WADDR[5], 1.0);
   $setup(posedge WADDR[6], posedge WCLKN, 1.0);
   $setup(negedge WADDR[6], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[6], 1.0);
   $hold(posedge WCLKN, negedge WADDR[6], 1.0);
   $setup(posedge WADDR[7], posedge WCLKN, 1.0);
   $setup(negedge WADDR[7], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[7], 1.0);
   $hold(posedge WCLKN, negedge WADDR[7], 1.0);
   $setup(posedge WADDR[8], posedge WCLKN, 1.0);
   $setup(negedge WADDR[8], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[8], 1.0);
   $hold(posedge WCLKN, negedge WADDR[8], 1.0);
   $setup(posedge WADDR[9], posedge WCLKN, 1.0);
   $setup(negedge WADDR[9], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[9], 1.0);
   $hold(posedge WCLKN, negedge WADDR[9], 1.0);
   $setup(posedge WADDR[10], posedge WCLKN, 1.0);
   $setup(negedge WADDR[10], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[10], 1.0);
   $hold(posedge WCLKN, negedge WADDR[10], 1.0);
   $setup(posedge WDATA[0], posedge WCLKN, 1.0);
   $setup(negedge WDATA[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[0], 1.0);
   $hold(posedge WCLKN, negedge WDATA[0], 1.0);
   $setup(posedge WDATA[1], posedge WCLKN, 1.0);
   $setup(negedge WDATA[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[1], 1.0);
   $hold(posedge WCLKN, negedge WDATA[1], 1.0);
   $setup(posedge WDATA[2], posedge WCLKN, 1.0);
   $setup(negedge WDATA[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[2], 1.0);
   $hold(posedge WCLKN, negedge WDATA[2], 1.0);
   $setup(posedge WDATA[3], posedge WCLKN, 1.0);
   $setup(negedge WDATA[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[3], 1.0);
   $hold(posedge WCLKN, negedge WDATA[3], 1.0);
   $setup(posedge WDATA[4], posedge WCLKN, 1.0);
   $setup(negedge WDATA[4], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[4], 1.0);
   $hold(posedge WCLKN, negedge WDATA[4], 1.0);
   $setup(posedge WDATA[5], posedge WCLKN, 1.0);
   $setup(negedge WDATA[5], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[5], 1.0);
   $hold(posedge WCLKN, negedge WDATA[5], 1.0);
   $setup(posedge WDATA[6], posedge WCLKN, 1.0);
   $setup(negedge WDATA[6], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[6], 1.0);
   $hold(posedge WCLKN, negedge WDATA[6], 1.0);
   $setup(posedge WDATA[7], posedge WCLKN, 1.0);
   $setup(negedge WDATA[7], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[7], 1.0);
   $hold(posedge WCLKN, negedge WDATA[7], 1.0);
   $setup(posedge WDATA[8], posedge WCLKN, 1.0);
   $setup(negedge WDATA[8], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[8], 1.0);
   $hold(posedge WCLKN, negedge WDATA[8], 1.0);
   $setup(posedge WDATA[9], posedge WCLKN, 1.0);
   $setup(negedge WDATA[9], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[9], 1.0);
   $hold(posedge WCLKN, negedge WDATA[9], 1.0);
   $setup(posedge WDATA[10], posedge WCLKN, 1.0);
   $setup(negedge WDATA[10], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[10], 1.0);
   $hold(posedge WCLKN, negedge WDATA[10], 1.0);
   $setup(posedge WDATA[11], posedge WCLKN, 1.0);
   $setup(negedge WDATA[11], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[11], 1.0);
   $hold(posedge WCLKN, negedge WDATA[11], 1.0);
   $setup(posedge WDATA[12], posedge WCLKN, 1.0);
   $setup(negedge WDATA[12], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[12], 1.0);
   $hold(posedge WCLKN, negedge WDATA[12], 1.0);
   $setup(posedge WDATA[13], posedge WCLKN, 1.0);
   $setup(negedge WDATA[13], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[13], 1.0);
   $hold(posedge WCLKN, negedge WDATA[13], 1.0);
   $setup(posedge WDATA[14], posedge WCLKN, 1.0);
   $setup(negedge WDATA[14], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[14], 1.0);
   $hold(posedge WCLKN, negedge WDATA[14], 1.0);
   $setup(posedge WDATA[15], posedge WCLKN, 1.0);
   $setup(negedge WDATA[15], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[15], 1.0);
   $hold(posedge WCLKN, negedge WDATA[15], 1.0);
   $setup(posedge WCLKE, posedge WCLKN, 1.0);
   $setup(negedge WCLKE, posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WCLKE, 1.0);
   $hold(posedge WCLKN, negedge WCLKE, 1.0);
   $setup(posedge WE, posedge WCLKN, 1.0);
   $setup(negedge WE, posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WE, 1.0);
   $hold(posedge WCLKN, negedge WE, 1.0);
   $setup(posedge RADDR[0], posedge RCLK, 1.0);
   $setup(negedge RADDR[0], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[0], 1.0);
   $hold(posedge RCLK, negedge RADDR[0], 1.0);
   $setup(posedge RADDR[1], posedge RCLK, 1.0);
   $setup(negedge RADDR[1], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[1], 1.0);
   $hold(posedge RCLK, negedge RADDR[1], 1.0);
   $setup(posedge RADDR[2], posedge RCLK, 1.0);
   $setup(negedge RADDR[2], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[2], 1.0);
   $hold(posedge RCLK, negedge RADDR[2], 1.0);
   $setup(posedge RADDR[3], posedge RCLK, 1.0);
   $setup(negedge RADDR[3], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[3], 1.0);
   $hold(posedge RCLK, negedge RADDR[3], 1.0);
   $setup(posedge RADDR[4], posedge RCLK, 1.0);
   $setup(negedge RADDR[4], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[4], 1.0);
   $hold(posedge RCLK, negedge RADDR[4], 1.0);
   $setup(posedge RADDR[5], posedge RCLK, 1.0);
   $setup(negedge RADDR[5], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[5], 1.0);
   $hold(posedge RCLK, negedge RADDR[5], 1.0);
   $setup(posedge RADDR[6], posedge RCLK, 1.0);
   $setup(negedge RADDR[6], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[6], 1.0);
   $hold(posedge RCLK, negedge RADDR[6], 1.0);
   $setup(posedge RADDR[7], posedge RCLK, 1.0);
   $setup(negedge RADDR[7], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[7], 1.0);
   $hold(posedge RCLK, negedge RADDR[7], 1.0);
   $setup(posedge RADDR[8], posedge RCLK, 1.0);
   $setup(negedge RADDR[8], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[8], 1.0);
   $hold(posedge RCLK, negedge RADDR[8], 1.0);
   $setup(posedge RADDR[9], posedge RCLK, 1.0);
   $setup(negedge RADDR[9], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[9], 1.0);
   $hold(posedge RCLK, negedge RADDR[9], 1.0);
   $setup(posedge RADDR[10], posedge RCLK, 1.0);
   $setup(negedge RADDR[10], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[10], 1.0);
   $hold(posedge RCLK, negedge RADDR[10], 1.0);
   $setup(posedge RCLKE, posedge RCLK, 1.0);
   $setup(negedge RCLKE, posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RCLKE, 1.0);
   $hold(posedge RCLK, negedge RCLKE, 1.0);
   $setup(posedge RE, posedge RCLK, 1.0);
   $setup(negedge RE, posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RE, 1.0);
   $hold(posedge RCLK, negedge RE, 1.0);

endspecify
`endif

endmodule //SB_RAM40_4KNW

`timescale 1ps/1ps
module SB_RAM40_4KNRNW (RDATA, RCLKN, RCLKE, RE, RADDR, WCLKN, WCLKE, WE, WADDR, MASK, WDATA);
output [15:0] RDATA;
input RCLKN;
input RCLKE;
input RE;
input [10:0] RADDR;
input WCLKN;
input WCLKE;
input WE;
input [10:0] WADDR;
input [15:0] MASK;
input [15:0] WDATA;

parameter WRITE_MODE = 0; /// can be integer 0(256X16 mode) or 1(512X8 mode) or 2(1024X4 mode) or 3(2048X2 mode)
parameter READ_MODE = 0;  /// can be integer 0(256X16 mode) or 1(512X8 mode) or 2(1024X4 mode) or 3(2048X2 mode)


parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

wire WCLK;
wire RCLK;
assign (weak0, weak1) RCLKE =1'b1 ;
assign (weak0, weak1) RE =1'b0 ;
assign (weak0, weak1) WCLKE =1'b1 ;
assign (weak0, weak1) WE =1'b0 ;
assign WCLK = ~WCLKN;
assign RCLK = ~RCLKN;

SB_RAM40_4K ram40_4K_nrnw_inst (
	.RDATA(RDATA),
	.RCLK(RCLK),
	.RCLKE(RCLKE),
	.RE(RE),
	.RADDR(RADDR),
	.WCLK(WCLK),
	.WCLKE(WCLKE),
	.WE(WE),
	.WADDR(WADDR),
	.MASK(MASK),
	.WDATA(WDATA));

defparam ram40_4K_nrnw_inst.WRITE_MODE = WRITE_MODE;
defparam ram40_4K_nrnw_inst.READ_MODE = READ_MODE;
defparam ram40_4K_nrnw_inst.INIT_0 = INIT_0;
defparam ram40_4K_nrnw_inst.INIT_1 = INIT_1;
defparam ram40_4K_nrnw_inst.INIT_2 = INIT_2;
defparam ram40_4K_nrnw_inst.INIT_3 = INIT_3;
defparam ram40_4K_nrnw_inst.INIT_4 = INIT_4;
defparam ram40_4K_nrnw_inst.INIT_5 = INIT_5;
defparam ram40_4K_nrnw_inst.INIT_6 = INIT_6;
defparam ram40_4K_nrnw_inst.INIT_7 = INIT_7;
defparam ram40_4K_nrnw_inst.INIT_8 = INIT_8;
defparam ram40_4K_nrnw_inst.INIT_9 = INIT_9;
defparam ram40_4K_nrnw_inst.INIT_A = INIT_A;
defparam ram40_4K_nrnw_inst.INIT_B = INIT_B;
defparam ram40_4K_nrnw_inst.INIT_C = INIT_C;
defparam ram40_4K_nrnw_inst.INIT_D = INIT_D;
defparam ram40_4K_nrnw_inst.INIT_E = INIT_E;
defparam ram40_4K_nrnw_inst.INIT_F = INIT_F;


`ifdef TIMINGCHECK
specify
   (RCLKN *> RDATA[0]) = (1.0, 1.0);
   (RCLKN *> RDATA[1]) = (1.0, 1.0);
   (RCLKN *> RDATA[2]) = (1.0, 1.0);
   (RCLKN *> RDATA[3]) = (1.0, 1.0);
   (RCLKN *> RDATA[4]) = (1.0, 1.0);
   (RCLKN *> RDATA[5]) = (1.0, 1.0);
   (RCLKN *> RDATA[6]) = (1.0, 1.0);
   (RCLKN *> RDATA[7]) = (1.0, 1.0);
   (RCLKN *> RDATA[8]) = (1.0, 1.0);
   (RCLKN *> RDATA[9]) = (1.0, 1.0);
   (RCLKN *> RDATA[10]) = (1.0, 1.0);
   (RCLKN *> RDATA[11]) = (1.0, 1.0);
   (RCLKN *> RDATA[12]) = (1.0, 1.0);
   (RCLKN *> RDATA[13]) = (1.0, 1.0);
   (RCLKN *> RDATA[14]) = (1.0, 1.0);
   (RCLKN *> RDATA[15]) = (1.0, 1.0);
   $setup(posedge MASK[0], posedge WCLKN, 1.0);
   $setup(negedge MASK[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[0], 1.0);
   $hold(posedge WCLKN, negedge MASK[0], 1.0);
   $setup(posedge MASK[1], posedge WCLKN, 1.0);
   $setup(negedge MASK[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[1], 1.0);
   $hold(posedge WCLKN, negedge MASK[1], 1.0);
   $setup(posedge MASK[2], posedge WCLKN, 1.0);
   $setup(negedge MASK[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[2], 1.0);
   $hold(posedge WCLKN, negedge MASK[2], 1.0);
   $setup(posedge MASK[3], posedge WCLKN, 1.0);
   $setup(negedge MASK[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[3], 1.0);
   $hold(posedge WCLKN, negedge MASK[3], 1.0);
   $setup(posedge MASK[4], posedge WCLKN, 1.0);
   $setup(negedge MASK[4], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[4], 1.0);
   $hold(posedge WCLKN, negedge MASK[4], 1.0);
   $setup(posedge MASK[5], posedge WCLKN, 1.0);
   $setup(negedge MASK[5], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[5], 1.0);
   $hold(posedge WCLKN, negedge MASK[5], 1.0);
   $setup(posedge MASK[6], posedge WCLKN, 1.0);
   $setup(negedge MASK[6], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[6], 1.0);
   $hold(posedge WCLKN, negedge MASK[6], 1.0);
   $setup(posedge MASK[7], posedge WCLKN, 1.0);
   $setup(negedge MASK[7], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[7], 1.0);
   $hold(posedge WCLKN, negedge MASK[7], 1.0);
   $setup(posedge MASK[8], posedge WCLKN, 1.0);
   $setup(negedge MASK[8], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[8], 1.0);
   $hold(posedge WCLKN, negedge MASK[8], 1.0);
   $setup(posedge MASK[9], posedge WCLKN, 1.0);
   $setup(negedge MASK[9], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[9], 1.0);
   $hold(posedge WCLKN, negedge MASK[9], 1.0);
   $setup(posedge MASK[10], posedge WCLKN, 1.0);
   $setup(negedge MASK[10], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[10], 1.0);
   $hold(posedge WCLKN, negedge MASK[10], 1.0);
   $setup(posedge MASK[11], posedge WCLKN, 1.0);
   $setup(negedge MASK[11], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[11], 1.0);
   $hold(posedge WCLKN, negedge MASK[11], 1.0);
   $setup(posedge MASK[12], posedge WCLKN, 1.0);
   $setup(negedge MASK[12], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[12], 1.0);
   $hold(posedge WCLKN, negedge MASK[12], 1.0);
   $setup(posedge MASK[13], posedge WCLKN, 1.0);
   $setup(negedge MASK[13], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[13], 1.0);
   $hold(posedge WCLKN, negedge MASK[13], 1.0);
   $setup(posedge MASK[14], posedge WCLKN, 1.0);
   $setup(negedge MASK[14], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[14], 1.0);
   $hold(posedge WCLKN, negedge MASK[14], 1.0);
   $setup(posedge MASK[15], posedge WCLKN, 1.0);
   $setup(negedge MASK[15], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[15], 1.0);
   $hold(posedge WCLKN, negedge MASK[15], 1.0);
   $setup(posedge WADDR[0], posedge WCLKN, 1.0);
   $setup(negedge WADDR[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[0], 1.0);
   $hold(posedge WCLKN, negedge WADDR[0], 1.0);
   $setup(posedge WADDR[1], posedge WCLKN, 1.0);
   $setup(negedge WADDR[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[1], 1.0);
   $hold(posedge WCLKN, negedge WADDR[1], 1.0);
   $setup(posedge WADDR[2], posedge WCLKN, 1.0);
   $setup(negedge WADDR[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[2], 1.0);
   $hold(posedge WCLKN, negedge WADDR[2], 1.0);
   $setup(posedge WADDR[3], posedge WCLKN, 1.0);
   $setup(negedge WADDR[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[3], 1.0);
   $hold(posedge WCLKN, negedge WADDR[3], 1.0);
   $setup(posedge WADDR[4], posedge WCLKN, 1.0);
   $setup(negedge WADDR[4], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[4], 1.0);
   $hold(posedge WCLKN, negedge WADDR[4], 1.0);
   $setup(posedge WADDR[5], posedge WCLKN, 1.0);
   $setup(negedge WADDR[5], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[5], 1.0);
   $hold(posedge WCLKN, negedge WADDR[5], 1.0);
   $setup(posedge WADDR[6], posedge WCLKN, 1.0);
   $setup(negedge WADDR[6], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[6], 1.0);
   $hold(posedge WCLKN, negedge WADDR[6], 1.0);
   $setup(posedge WADDR[7], posedge WCLKN, 1.0);
   $setup(negedge WADDR[7], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[7], 1.0);
   $hold(posedge WCLKN, negedge WADDR[7], 1.0);
   $setup(posedge WADDR[8], posedge WCLKN, 1.0);
   $setup(negedge WADDR[8], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[8], 1.0);
   $hold(posedge WCLKN, negedge WADDR[8], 1.0);
   $setup(posedge WADDR[9], posedge WCLKN, 1.0);
   $setup(negedge WADDR[9], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[9], 1.0);
   $hold(posedge WCLKN, negedge WADDR[9], 1.0);
   $setup(posedge WADDR[10], posedge WCLKN, 1.0);
   $setup(negedge WADDR[10], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[10], 1.0);
   $hold(posedge WCLKN, negedge WADDR[10], 1.0);
   $setup(posedge WDATA[0], posedge WCLKN, 1.0);
   $setup(negedge WDATA[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[0], 1.0);
   $hold(posedge WCLKN, negedge WDATA[0], 1.0);
   $setup(posedge WDATA[1], posedge WCLKN, 1.0);
   $setup(negedge WDATA[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[1], 1.0);
   $hold(posedge WCLKN, negedge WDATA[1], 1.0);
   $setup(posedge WDATA[2], posedge WCLKN, 1.0);
   $setup(negedge WDATA[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[2], 1.0);
   $hold(posedge WCLKN, negedge WDATA[2], 1.0);
   $setup(posedge WDATA[3], posedge WCLKN, 1.0);
   $setup(negedge WDATA[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[3], 1.0);
   $hold(posedge WCLKN, negedge WDATA[3], 1.0);
   $setup(posedge WDATA[4], posedge WCLKN, 1.0);
   $setup(negedge WDATA[4], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[4], 1.0);
   $hold(posedge WCLKN, negedge WDATA[4], 1.0);
   $setup(posedge WDATA[5], posedge WCLKN, 1.0);
   $setup(negedge WDATA[5], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[5], 1.0);
   $hold(posedge WCLKN, negedge WDATA[5], 1.0);
   $setup(posedge WDATA[6], posedge WCLKN, 1.0);
   $setup(negedge WDATA[6], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[6], 1.0);
   $hold(posedge WCLKN, negedge WDATA[6], 1.0);
   $setup(posedge WDATA[7], posedge WCLKN, 1.0);
   $setup(negedge WDATA[7], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[7], 1.0);
   $hold(posedge WCLKN, negedge WDATA[7], 1.0);
   $setup(posedge WDATA[8], posedge WCLKN, 1.0);
   $setup(negedge WDATA[8], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[8], 1.0);
   $hold(posedge WCLKN, negedge WDATA[8], 1.0);
   $setup(posedge WDATA[9], posedge WCLKN, 1.0);
   $setup(negedge WDATA[9], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[9], 1.0);
   $hold(posedge WCLKN, negedge WDATA[9], 1.0);
   $setup(posedge WDATA[10], posedge WCLKN, 1.0);
   $setup(negedge WDATA[10], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[10], 1.0);
   $hold(posedge WCLKN, negedge WDATA[10], 1.0);
   $setup(posedge WDATA[11], posedge WCLKN, 1.0);
   $setup(negedge WDATA[11], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[11], 1.0);
   $hold(posedge WCLKN, negedge WDATA[11], 1.0);
   $setup(posedge WDATA[12], posedge WCLKN, 1.0);
   $setup(negedge WDATA[12], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[12], 1.0);
   $hold(posedge WCLKN, negedge WDATA[12], 1.0);
   $setup(posedge WDATA[13], posedge WCLKN, 1.0);
   $setup(negedge WDATA[13], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[13], 1.0);
   $hold(posedge WCLKN, negedge WDATA[13], 1.0);
   $setup(posedge WDATA[14], posedge WCLKN, 1.0);
   $setup(negedge WDATA[14], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[14], 1.0);
   $hold(posedge WCLKN, negedge WDATA[14], 1.0);
   $setup(posedge WDATA[15], posedge WCLKN, 1.0);
   $setup(negedge WDATA[15], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[15], 1.0);
   $hold(posedge WCLKN, negedge WDATA[15], 1.0);
   $setup(posedge WCLKE, posedge WCLKN, 1.0);
   $setup(negedge WCLKE, posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WCLKE, 1.0);
   $hold(posedge WCLKN, negedge WCLKE, 1.0);
   $setup(posedge WE, posedge WCLKN, 1.0);
   $setup(negedge WE, posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WE, 1.0);
   $hold(posedge WCLKN, negedge WE, 1.0);
   $setup(posedge RADDR[0], posedge RCLKN, 1.0);
   $setup(negedge RADDR[0], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[0], 1.0);
   $hold(posedge RCLKN, negedge RADDR[0], 1.0);
   $setup(posedge RADDR[1], posedge RCLKN, 1.0);
   $setup(negedge RADDR[1], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[1], 1.0);
   $hold(posedge RCLKN, negedge RADDR[1], 1.0);
   $setup(posedge RADDR[2], posedge RCLKN, 1.0);
   $setup(negedge RADDR[2], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[2], 1.0);
   $hold(posedge RCLKN, negedge RADDR[2], 1.0);
   $setup(posedge RADDR[3], posedge RCLKN, 1.0);
   $setup(negedge RADDR[3], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[3], 1.0);
   $hold(posedge RCLKN, negedge RADDR[3], 1.0);
   $setup(posedge RADDR[4], posedge RCLKN, 1.0);
   $setup(negedge RADDR[4], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[4], 1.0);
   $hold(posedge RCLKN, negedge RADDR[4], 1.0);
   $setup(posedge RADDR[5], posedge RCLKN, 1.0);
   $setup(negedge RADDR[5], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[5], 1.0);
   $hold(posedge RCLKN, negedge RADDR[5], 1.0);
   $setup(posedge RADDR[6], posedge RCLKN, 1.0);
   $setup(negedge RADDR[6], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[6], 1.0);
   $hold(posedge RCLKN, negedge RADDR[6], 1.0);
   $setup(posedge RADDR[7], posedge RCLKN, 1.0);
   $setup(negedge RADDR[7], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[7], 1.0);
   $hold(posedge RCLKN, negedge RADDR[7], 1.0);
   $setup(posedge RADDR[8], posedge RCLKN, 1.0);
   $setup(negedge RADDR[8], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[8], 1.0);
   $hold(posedge RCLKN, negedge RADDR[8], 1.0);
   $setup(posedge RADDR[9], posedge RCLKN, 1.0);
   $setup(negedge RADDR[9], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[9], 1.0);
   $hold(posedge RCLKN, negedge RADDR[9], 1.0);
   $setup(posedge RADDR[10], posedge RCLKN, 1.0);
   $setup(negedge RADDR[10], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[10], 1.0);
   $hold(posedge RCLKN, negedge RADDR[10], 1.0);
   $setup(posedge RCLKE, posedge RCLKN, 1.0);
   $setup(negedge RCLKE, posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RCLKE, 1.0);
   $hold(posedge RCLKN, negedge RCLKE, 1.0);
   $setup(posedge RE, posedge RCLKN, 1.0);
   $setup(negedge RE, posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RE, 1.0);
   $hold(posedge RCLKN, negedge RE, 1.0);

endspecify
`endif

endmodule //SB_RAM40_4KNRNW

`timescale 1ps/1ps
module SB_RAM40_4K (RDATA, RCLK, RCLKE, RE, RADDR, WCLK, WCLKE, WE, WADDR, MASK, WDATA);
output [15:0] RDATA;
input RCLK;
input RCLKE;
input RE;
input [10:0] RADDR;
input WCLK;
input WCLKE;
input WE;
input [10:0] WADDR;
input [15:0] MASK;
input [15:0] WDATA;

assign (weak0, weak1) MASK = 16'b0;

parameter WRITE_MODE = 0; /// can be integer 0(256X16 mode) or 1(512X8 mode) or 2(1024X4 mode) or 3(2048X2 mode)
parameter READ_MODE = 0;  /// can be integer 0(256X16 mode) or 1(512X8 mode) or 2(1024X4 mode) or 3(2048X2 mode)


parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

wire [15:0] RD;
wire [15:0] WD;
wire [15:0] MASK_RAM;

reg [10:8] RADDR_reg;
always @(posedge RCLK) begin
	RADDR_reg[10:8] <= RADDR[10:8];
end

read_data_decoder read_decoder_inst (
	.di(RD),
	.ai(RADDR_reg[10:8]),
	.do(RDATA)
);
defparam read_decoder_inst.READ_MODE = READ_MODE;

write_data_decoder write_decoder_inst (
	.di(WDATA),
	.do(WD)
);
defparam write_decoder_inst.WRITE_MODE = WRITE_MODE;

mask_decoder mask_decoder_inst(
	.mi(MASK),
	.ai(WADDR[10:8]),
	.mo(MASK_RAM)
);
defparam mask_decoder_inst.WRITE_MODE = WRITE_MODE;

SB_RAM4K ram_inst (
	.RDATA(RD),
	.RCLK(RCLK),
	.RCLKE(RCLKE),
	.RE(RE),
	.RADDR(RADDR[7:0]),
	.WCLK(WCLK),
	.WCLKE(WCLKE),
	.WE(WE),
	.WADDR(WADDR[7:0]),
	.MASK(MASK_RAM),
	.WDATA(WD));

defparam ram_inst.INIT_0 = INIT_0;
defparam ram_inst.INIT_1 = INIT_1;
defparam ram_inst.INIT_2 = INIT_2;
defparam ram_inst.INIT_3 = INIT_3;
defparam ram_inst.INIT_4 = INIT_4;
defparam ram_inst.INIT_5 = INIT_5;
defparam ram_inst.INIT_6 = INIT_6;
defparam ram_inst.INIT_7 = INIT_7;
defparam ram_inst.INIT_8 = INIT_8;
defparam ram_inst.INIT_9 = INIT_9;
defparam ram_inst.INIT_A = INIT_A;
defparam ram_inst.INIT_B = INIT_B;
defparam ram_inst.INIT_C = INIT_C;
defparam ram_inst.INIT_D = INIT_D;
defparam ram_inst.INIT_E = INIT_E;
defparam ram_inst.INIT_F = INIT_F;

`ifdef TIMINGCHECK
specify
   (RCLK *> RDATA[0]) = (1.0, 1.0);
   (RCLK *> RDATA[1]) = (1.0, 1.0);
   (RCLK *> RDATA[2]) = (1.0, 1.0);
   (RCLK *> RDATA[3]) = (1.0, 1.0);
   (RCLK *> RDATA[4]) = (1.0, 1.0);
   (RCLK *> RDATA[5]) = (1.0, 1.0);
   (RCLK *> RDATA[6]) = (1.0, 1.0);
   (RCLK *> RDATA[7]) = (1.0, 1.0);
   (RCLK *> RDATA[8]) = (1.0, 1.0);
   (RCLK *> RDATA[9]) = (1.0, 1.0);
   (RCLK *> RDATA[10]) = (1.0, 1.0);
   (RCLK *> RDATA[11]) = (1.0, 1.0);
   (RCLK *> RDATA[12]) = (1.0, 1.0);
   (RCLK *> RDATA[13]) = (1.0, 1.0);
   (RCLK *> RDATA[14]) = (1.0, 1.0);
   (RCLK *> RDATA[15]) = (1.0, 1.0);
   $setup(posedge MASK[0], posedge WCLK, 1.0);
   $setup(negedge MASK[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[0], 1.0);
   $hold(posedge WCLK, negedge MASK[0], 1.0);
   $setup(posedge MASK[1], posedge WCLK, 1.0);
   $setup(negedge MASK[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[1], 1.0);
   $hold(posedge WCLK, negedge MASK[1], 1.0);
   $setup(posedge MASK[2], posedge WCLK, 1.0);
   $setup(negedge MASK[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[2], 1.0);
   $hold(posedge WCLK, negedge MASK[2], 1.0);
   $setup(posedge MASK[3], posedge WCLK, 1.0);
   $setup(negedge MASK[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[3], 1.0);
   $hold(posedge WCLK, negedge MASK[3], 1.0);
   $setup(posedge MASK[4], posedge WCLK, 1.0);
   $setup(negedge MASK[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[4], 1.0);
   $hold(posedge WCLK, negedge MASK[4], 1.0);
   $setup(posedge MASK[5], posedge WCLK, 1.0);
   $setup(negedge MASK[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[5], 1.0);
   $hold(posedge WCLK, negedge MASK[5], 1.0);
   $setup(posedge MASK[6], posedge WCLK, 1.0);
   $setup(negedge MASK[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[6], 1.0);
   $hold(posedge WCLK, negedge MASK[6], 1.0);
   $setup(posedge MASK[7], posedge WCLK, 1.0);
   $setup(negedge MASK[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[7], 1.0);
   $hold(posedge WCLK, negedge MASK[7], 1.0);
   $setup(posedge MASK[8], posedge WCLK, 1.0);
   $setup(negedge MASK[8], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[8], 1.0);
   $hold(posedge WCLK, negedge MASK[8], 1.0);
   $setup(posedge MASK[9], posedge WCLK, 1.0);
   $setup(negedge MASK[9], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[9], 1.0);
   $hold(posedge WCLK, negedge MASK[9], 1.0);
   $setup(posedge MASK[10], posedge WCLK, 1.0);
   $setup(negedge MASK[10], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[10], 1.0);
   $hold(posedge WCLK, negedge MASK[10], 1.0);
   $setup(posedge MASK[11], posedge WCLK, 1.0);
   $setup(negedge MASK[11], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[11], 1.0);
   $hold(posedge WCLK, negedge MASK[11], 1.0);
   $setup(posedge MASK[12], posedge WCLK, 1.0);
   $setup(negedge MASK[12], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[12], 1.0);
   $hold(posedge WCLK, negedge MASK[12], 1.0);
   $setup(posedge MASK[13], posedge WCLK, 1.0);
   $setup(negedge MASK[13], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[13], 1.0);
   $hold(posedge WCLK, negedge MASK[13], 1.0);
   $setup(posedge MASK[14], posedge WCLK, 1.0);
   $setup(negedge MASK[14], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[14], 1.0);
   $hold(posedge WCLK, negedge MASK[14], 1.0);
   $setup(posedge MASK[15], posedge WCLK, 1.0);
   $setup(negedge MASK[15], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[15], 1.0);
   $hold(posedge WCLK, negedge MASK[15], 1.0);
   $setup(posedge WADDR[0], posedge WCLK, 1.0);
   $setup(negedge WADDR[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[0], 1.0);
   $hold(posedge WCLK, negedge WADDR[0], 1.0);
   $setup(posedge WADDR[1], posedge WCLK, 1.0);
   $setup(negedge WADDR[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[1], 1.0);
   $hold(posedge WCLK, negedge WADDR[1], 1.0);
   $setup(posedge WADDR[2], posedge WCLK, 1.0);
   $setup(negedge WADDR[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[2], 1.0);
   $hold(posedge WCLK, negedge WADDR[2], 1.0);
   $setup(posedge WADDR[3], posedge WCLK, 1.0);
   $setup(negedge WADDR[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[3], 1.0);
   $hold(posedge WCLK, negedge WADDR[3], 1.0);
   $setup(posedge WADDR[4], posedge WCLK, 1.0);
   $setup(negedge WADDR[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[4], 1.0);
   $hold(posedge WCLK, negedge WADDR[4], 1.0);
   $setup(posedge WADDR[5], posedge WCLK, 1.0);
   $setup(negedge WADDR[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[5], 1.0);
   $hold(posedge WCLK, negedge WADDR[5], 1.0);
   $setup(posedge WADDR[6], posedge WCLK, 1.0);
   $setup(negedge WADDR[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[6], 1.0);
   $hold(posedge WCLK, negedge WADDR[6], 1.0);
   $setup(posedge WADDR[7], posedge WCLK, 1.0);
   $setup(negedge WADDR[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[7], 1.0);
   $hold(posedge WCLK, negedge WADDR[7], 1.0);
   $setup(posedge WADDR[8], posedge WCLK, 1.0);
   $setup(negedge WADDR[8], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[8], 1.0);
   $hold(posedge WCLK, negedge WADDR[8], 1.0);
   $setup(posedge WADDR[9], posedge WCLK, 1.0);
   $setup(negedge WADDR[9], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[9], 1.0);
   $hold(posedge WCLK, negedge WADDR[9], 1.0);
   $setup(posedge WADDR[10], posedge WCLK, 1.0);
   $setup(negedge WADDR[10], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[10], 1.0);
   $hold(posedge WCLK, negedge WADDR[10], 1.0);
   $setup(posedge WDATA[0], posedge WCLK, 1.0);
   $setup(negedge WDATA[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[0], 1.0);
   $hold(posedge WCLK, negedge WDATA[0], 1.0);
   $setup(posedge WDATA[1], posedge WCLK, 1.0);
   $setup(negedge WDATA[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[1], 1.0);
   $hold(posedge WCLK, negedge WDATA[1], 1.0);
   $setup(posedge WDATA[2], posedge WCLK, 1.0);
   $setup(negedge WDATA[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[2], 1.0);
   $hold(posedge WCLK, negedge WDATA[2], 1.0);
   $setup(posedge WDATA[3], posedge WCLK, 1.0);
   $setup(negedge WDATA[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[3], 1.0);
   $hold(posedge WCLK, negedge WDATA[3], 1.0);
   $setup(posedge WDATA[4], posedge WCLK, 1.0);
   $setup(negedge WDATA[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[4], 1.0);
   $hold(posedge WCLK, negedge WDATA[4], 1.0);
   $setup(posedge WDATA[5], posedge WCLK, 1.0);
   $setup(negedge WDATA[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[5], 1.0);
   $hold(posedge WCLK, negedge WDATA[5], 1.0);
   $setup(posedge WDATA[6], posedge WCLK, 1.0);
   $setup(negedge WDATA[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[6], 1.0);
   $hold(posedge WCLK, negedge WDATA[6], 1.0);
   $setup(posedge WDATA[7], posedge WCLK, 1.0);
   $setup(negedge WDATA[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[7], 1.0);
   $hold(posedge WCLK, negedge WDATA[7], 1.0);
   $setup(posedge WDATA[8], posedge WCLK, 1.0);
   $setup(negedge WDATA[8], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[8], 1.0);
   $hold(posedge WCLK, negedge WDATA[8], 1.0);
   $setup(posedge WDATA[9], posedge WCLK, 1.0);
   $setup(negedge WDATA[9], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[9], 1.0);
   $hold(posedge WCLK, negedge WDATA[9], 1.0);
   $setup(posedge WDATA[10], posedge WCLK, 1.0);
   $setup(negedge WDATA[10], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[10], 1.0);
   $hold(posedge WCLK, negedge WDATA[10], 1.0);
   $setup(posedge WDATA[11], posedge WCLK, 1.0);
   $setup(negedge WDATA[11], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[11], 1.0);
   $hold(posedge WCLK, negedge WDATA[11], 1.0);
   $setup(posedge WDATA[12], posedge WCLK, 1.0);
   $setup(negedge WDATA[12], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[12], 1.0);
   $hold(posedge WCLK, negedge WDATA[12], 1.0);
   $setup(posedge WDATA[13], posedge WCLK, 1.0);
   $setup(negedge WDATA[13], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[13], 1.0);
   $hold(posedge WCLK, negedge WDATA[13], 1.0);
   $setup(posedge WDATA[14], posedge WCLK, 1.0);
   $setup(negedge WDATA[14], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[14], 1.0);
   $hold(posedge WCLK, negedge WDATA[14], 1.0);
   $setup(posedge WDATA[15], posedge WCLK, 1.0);
   $setup(negedge WDATA[15], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[15], 1.0);
   $hold(posedge WCLK, negedge WDATA[15], 1.0);
   $setup(posedge WCLKE, posedge WCLK, 1.0);
   $setup(negedge WCLKE, posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WCLKE, 1.0);
   $hold(posedge WCLK, negedge WCLKE, 1.0);
   $setup(posedge WE, posedge WCLK, 1.0);
   $setup(negedge WE, posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WE, 1.0);
   $hold(posedge WCLK, negedge WE, 1.0);
   $setup(posedge RADDR[0], posedge RCLK, 1.0);
   $setup(negedge RADDR[0], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[0], 1.0);
   $hold(posedge RCLK, negedge RADDR[0], 1.0);
   $setup(posedge RADDR[1], posedge RCLK, 1.0);
   $setup(negedge RADDR[1], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[1], 1.0);
   $hold(posedge RCLK, negedge RADDR[1], 1.0);
   $setup(posedge RADDR[2], posedge RCLK, 1.0);
   $setup(negedge RADDR[2], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[2], 1.0);
   $hold(posedge RCLK, negedge RADDR[2], 1.0);
   $setup(posedge RADDR[3], posedge RCLK, 1.0);
   $setup(negedge RADDR[3], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[3], 1.0);
   $hold(posedge RCLK, negedge RADDR[3], 1.0);
   $setup(posedge RADDR[4], posedge RCLK, 1.0);
   $setup(negedge RADDR[4], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[4], 1.0);
   $hold(posedge RCLK, negedge RADDR[4], 1.0);
   $setup(posedge RADDR[5], posedge RCLK, 1.0);
   $setup(negedge RADDR[5], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[5], 1.0);
   $hold(posedge RCLK, negedge RADDR[5], 1.0);
   $setup(posedge RADDR[6], posedge RCLK, 1.0);
   $setup(negedge RADDR[6], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[6], 1.0);
   $hold(posedge RCLK, negedge RADDR[6], 1.0);
   $setup(posedge RADDR[7], posedge RCLK, 1.0);
   $setup(negedge RADDR[7], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[7], 1.0);
   $hold(posedge RCLK, negedge RADDR[7], 1.0);
   $setup(posedge RADDR[8], posedge RCLK, 1.0);
   $setup(negedge RADDR[8], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[8], 1.0);
   $hold(posedge RCLK, negedge RADDR[8], 1.0);
   $setup(posedge RADDR[9], posedge RCLK, 1.0);
   $setup(negedge RADDR[9], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[9], 1.0);
   $hold(posedge RCLK, negedge RADDR[9], 1.0);
   $setup(posedge RADDR[10], posedge RCLK, 1.0);
   $setup(negedge RADDR[10], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[10], 1.0);
   $hold(posedge RCLK, negedge RADDR[10], 1.0);
   $setup(posedge RCLKE, posedge RCLK, 1.0);
   $setup(negedge RCLKE, posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RCLKE, 1.0);
   $hold(posedge RCLK, negedge RCLKE, 1.0);
   $setup(posedge RE, posedge RCLK, 1.0);
   $setup(negedge RE, posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RE, 1.0);
   $hold(posedge RCLK, negedge RE, 1.0);

endspecify
`endif

endmodule //SB_RAM40_4K

`timescale 1ps/1ps

module read_data_decoder (
	di,
	ai,
	do
);

parameter READ_MODE = 0;

input [15:0] di;
input [2:0] ai;
output [15:0] do;
reg [15:0] do;

reg [1:0]mode;

initial 
begin
	if(READ_MODE == 0)
		mode = 2'b00;
	else if(READ_MODE == 1)
		mode = 2'b01;
	else if(READ_MODE == 2)
		mode = 2'b10;
	else if(READ_MODE == 3)
		mode = 2'b11;
	else
	begin
		$display (" SBT ERROR :  Unknown RAM READ MODE\n");
		$display (" Valid Modes are : 0, 1, 2, 3\n");
		//$display (" 0 -- 256X16 mode \n 1-- 512X8 mode \n 2 -- 1024X4 mode \n 3 -- 2048X2  mode \n");
		$finish;
	end
end

always @(mode, di, ai)
begin
	casex({mode,ai})
		5'b00xxx: do = di;
		5'b01xx0: do = {1'b0,di[14],1'b0,di[12],1'b0,di[10],1'b0,di[8],1'b0,di[6],1'b0,di[4],1'b0,di[2],1'b0,di[0]};
		5'b01xx1: do = {1'b0,di[15],1'b0,di[13],1'b0,di[11],1'b0,di[9],1'b0,di[7],1'b0,di[5],1'b0,di[3],1'b0,di[1]};
		5'b10x00: do = {1'b0,1'b0,di[12],1'b0,1'b0,1'b0,di[8],1'b0,1'b0,1'b0,di[4],1'b0,1'b0,1'b0,di[0],1'b0};
		5'b10x01: do = {1'b0,1'b0,di[13],1'b0,1'b0,1'b0,di[9],1'b0,1'b0,1'b0,di[5],1'b0,1'b0,1'b0,di[1],1'b0};
		5'b10x10: do = {1'b0,1'b0,di[14],1'b0,1'b0,1'b0,di[10],1'b0,1'b0,1'b0,di[6],1'b0,1'b0,1'b0,di[2],1'b0};
		5'b10x11: do = {1'b0,1'b0,di[15],1'b0,1'b0,1'b0,di[11],1'b0,1'b0,1'b0,di[7],1'b0,1'b0,1'b0,di[3],1'b0};
		5'b11000: do = {1'b0,1'b0,1'b0,1'b0,di[8],1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,di[0],1'b0,1'b0,1'b0};
		5'b11001: do = {1'b0,1'b0,1'b0,1'b0,di[9],1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,di[1],1'b0,1'b0,1'b0};
		5'b11010: do = {1'b0,1'b0,1'b0,1'b0,di[10],1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,di[2],1'b0,1'b0,1'b0};
		5'b11011: do = {1'b0,1'b0,1'b0,1'b0,di[11],1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,di[3],1'b0,1'b0,1'b0};
		5'b11100: do = {1'b0,1'b0,1'b0,1'b0,di[12],1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,di[4],1'b0,1'b0,1'b0};
		5'b11101: do = {1'b0,1'b0,1'b0,1'b0,di[13],1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,di[5],1'b0,1'b0,1'b0};
		5'b11110: do = {1'b0,1'b0,1'b0,1'b0,di[14],1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,di[6],1'b0,1'b0,1'b0};
		5'b11111: do = {1'b0,1'b0,1'b0,1'b0,di[15],1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,di[7],1'b0,1'b0,1'b0};
		default:
		begin
			$display ("SBT ERROR: End up in unknown address\n");
			$finish;
		end
	endcase
end

endmodule  // read_data_decoder

`timescale 1ps/1ps
module write_data_decoder (
	di,
	do
);

parameter WRITE_MODE = 0;

input [15:0] di;
output [15:0] do;

reg [15:0] do;


reg [1:0]mode;

initial 
begin
	if(WRITE_MODE == 0)
		mode = 2'b00;
	else if(WRITE_MODE == 1)
		mode = 2'b01;
	else if(WRITE_MODE == 2)
		mode = 2'b10;
	else if(WRITE_MODE == 3)
		mode = 2'b11;
	else
	begin
		$display (" SBT ERROR :  Unknown RAM WRITE MODE\n");
		$display (" Valid Modes are : 0, 1, 2, 3\n");
		//$display (" 0 -- 256X16 mode \n 1-- 512X8 mode \n 2 -- 1024X4 mode \n 3 -- 2048X2  mode \n");
		$finish;
	end
end

always @(mode, di )
begin
	case(mode)
		2'b00: do = di;
		2'b01: do = {di[14],di[14],di[12],di[12],di[10],di[10],di[8],di[8],di[6],di[6],di[4],di[4],di[2],di[2],di[0],di[0]};
		2'b10: do = {di[13],di[13],di[13],di[13],di[9],di[9],di[9],di[9],di[5],di[5],di[5],di[5],di[1],di[1],di[1],di[1]};
		2'b11: do = {di[11],di[11],di[11],di[11],di[11],di[11],di[11],di[11],di[3],di[3],di[3],di[3],di[3],di[3],di[3],di[3]};
	endcase
end

endmodule  // write_data_decoder

`timescale 1ps/1ps
module mask_decoder (
	mi,
	ai,
	mo
);

parameter WRITE_MODE = 0;

input [15:0] mi;
input [2:0] ai;
output [15:0] mo;

reg [15:0] mo;

reg [1:0]mode;

initial 
begin
	if(WRITE_MODE == 0)
		mode = 2'b00;
	else if(WRITE_MODE == 1)
		mode = 2'b01;
	else if(WRITE_MODE == 2)
		mode = 2'b10;
	else if(WRITE_MODE == 3)
		mode = 2'b11;
	else
	begin
		$display (" SBT ERROR :  Unknown RAM WRITE MODE\n");
		$display (" Valid Modes are : 0, 1, 2, 3\n");
		//$display (" 0 -- 256X16 mode \n 1-- 512X8 mode \n 2 -- 1024X4 mode \n 3 -- 2048X2  mode \n");
		$finish;
	end
end

always @(mode, mi, ai )
begin
	casex({mode,ai})
		5'b00xxx: mo = mi;
		5'b01xx0: mo = 16'hAAAA;
		5'b01xx1: mo = 16'h5555;
		5'b10x00: mo = 16'hEEEE;
		5'b10x01: mo = 16'hDDDD;
		5'b10x10: mo = 16'hBBBB;
		5'b10x11: mo = 16'h7777;
		5'b11000: mo = 16'hFEFE;
		5'b11001: mo = 16'hFDFD;
		5'b11010: mo = 16'hFBFB;
		5'b11011: mo = 16'hF7F7;
		5'b11100: mo = 16'hEFEF;
		5'b11101: mo = 16'hDFDF;
		5'b11110: mo = 16'hBFBF;
		5'b11111: mo = 16'h7F7F;
		default : 
		begin
			$display ("SBT ERROR: End up in unknown address\n");
			$finish;
		end
	endcase
end

endmodule  // mask_decoder

`timescale 1ps/1ps
module SB_RAM256x16 (RDATA, RCLK, RCLKE, RE, RADDR, WCLK, WCLKE, WE, WADDR, MASK, WDATA);
output [15:0] RDATA;
input RCLK;
input RCLKE;
input RE;
input [7:0] RADDR;
input WCLK;
input WCLKE;
input WE;
input [7:0] WADDR;
input [15:0] MASK;
input [15:0] WDATA;

parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

// local Parameters
localparam			CLOCK_PERIOD = 200;	//
localparam 			DELAY	= (CLOCK_PERIOD/10);		// Clock-to-output delay. Zero
							// time delays can be confusing
							// and sometimes cause problems.
localparam 			BUS_WIDTH = 16;		// Width of RAM (number of bits)

localparam 			ADDRESS_BUS_SIZE = 8;	// Number of bits required to
							// represent the RAM address

localparam   ADDRESSABLE_SPACE  = 2**ADDRESS_BUS_SIZE;	// Decimal address range [2^Size:0]


// SIGNAL DECLARATIONS
wire			   	WCLK_g, RCLK_g;
reg 				WCLKE_sync, RCLKE_sync; 
assign (weak0, weak1) RCLKE =1'b1 ;
assign (weak0, weak1) RE =1'b0 ;
assign (weak0, weak1) WCLKE =1'b1 ;
assign (weak0, weak1) WE =1'b0 ;
reg	Memory	[BUS_WIDTH*ADDRESSABLE_SPACE-1:0];
// 
event Read_e, Write_e;

//////////////////// Collision detect begins here ///////////////////////////////
localparam 	TRUE = 1'b1;
localparam	FALSE = 1'b0;
reg 		Time_Collision_Detected = 1'b0;
wire		Address_Collision_Detected;

event Collision_e;

time COLLISION_TIME_WINDOW = (CLOCK_PERIOD/8); // This is an arbitray value, but is better than using an absolute 
						    // value, because the actual time window depends on the actual silicon 
						    // implementation. Thus the test is indicative of an Error and not
						    // guaranteed to be an error. Even so this is usefull.
time time_WCLK_RCLK, time_WCLK, time_RCLK;


//function reg Check_Timed_Window_Violation;
function	Check_Timed_Window_Violation;	
input T1, T2, Minimum_Time_Window;
time T1, T2;
time Minimum_Time_Window;
time Difference;	
	begin
		Difference = (T1 - T2);
		if (Difference < 0) Difference = -Difference;
		Check_Timed_Window_Violation = (Difference < Minimum_Time_Window);
	end
endfunction


initial begin
       time_WCLK = CLOCK_PERIOD;	// Arbitrary initialisation value, ensure no window collison error on first clock edge.
       time_RCLK = (CLOCK_PERIOD*8);	// Arbitrary initialisation difference value, ensure no collision error on first clock edge.					
end

integer	i,j;


initial	//	initialize ram_4k by parameter, section by section
begin
	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[BUS_WIDTH*i+j]	=	INIT_0[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*1+BUS_WIDTH*i+j]	=	INIT_1[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*2+BUS_WIDTH*i+j]	=	INIT_2[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*3+BUS_WIDTH*i+j]	=	INIT_3[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*4+BUS_WIDTH*i+j]	=	INIT_4[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*5+BUS_WIDTH*i+j]	=	INIT_5[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*6+BUS_WIDTH*i+j]	=	INIT_6[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*7+BUS_WIDTH*i+j]	=	INIT_7[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*8+BUS_WIDTH*i+j]	=	INIT_8[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*9+BUS_WIDTH*i+j]	=	INIT_9[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*10+BUS_WIDTH*i+j]	=	INIT_A[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*11+BUS_WIDTH*i+j]	=	INIT_B[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*12+BUS_WIDTH*i+j]	=	INIT_C[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*13+BUS_WIDTH*i+j]	=	INIT_D[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*14+BUS_WIDTH*i+j]	=	INIT_E[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*15+BUS_WIDTH*i+j]	=	INIT_F[BUS_WIDTH*i+j];
	end

end

assign Address_Collision_Detected = ((RE & WE & WCLKE & RCLKE)&(WADDR == RADDR)); 

always @(WCLK or WCLKE) 
begin 
	if(~WCLK)
	WCLKE_sync = WCLKE;   	
end 

always @(RCLK or RCLKE) 
begin 
	if (~RCLK)
	RCLKE_sync = RCLKE; 	
end 

assign WCLK_g = WCLK & WCLKE_sync;
assign RCLK_g = RCLK & RCLKE_sync;


always @(posedge WCLK_g) begin
	time_WCLK = $time;
end

always @(posedge RCLK_g) begin
    	time_RCLK = $time;
end
integer	SB_RAM256X16_RDATA_log_file;					//.....................
initial	SB_RAM256X16_RDATA_log_file=("SB_RAM256X16_RDATA_log_file.txt");	//.....................
always @(posedge WCLK_g) begin

	Time_Collision_Detected = Check_Timed_Window_Violation(time_WCLK,time_RCLK,COLLISION_TIME_WINDOW);
        if (Time_Collision_Detected & Address_Collision_Detected)begin
        	$display("Warning: Write-Read collision detected, Data read value is XXXX\n");
 		$display("WCLK Time: %.3f   RCLK Time:%.3f  ",time_WCLK, time_RCLK,"WADDR: %d   RADDR:%d\n",WADDR, RADDR); 
 		$fdisplay(SB_RAM256X16_RDATA_log_file,"Warning: Write-Read collision detected, Data read value is XXXX\n");
		$fdisplay(SB_RAM256X16_RDATA_log_file,"WCLK Time: %.3f   RCLK Time:%.3f  ",time_WCLK, time_RCLK, "WADDR: %d   RADDR:%d\n",WADDR, RADDR); 	
 		-> Collision_e;
	end
end




//	code modify for universal verilog compiler

always @ (posedge WCLK_g)
begin
	if	(WE)
	begin
		-> Write_e;
		for	(i=0;i<=BUS_WIDTH-1; i=i+1)
		begin
			if	(MASK[i] !=1)
				Memory[WADDR*BUS_WIDTH+i]	<=	WDATA[i];
			else
				Memory[WADDR*BUS_WIDTH+i]	<=	Memory[WADDR*BUS_WIDTH+i];
		end
	end
end

//reg	[15:0]	RDATA = 0;
reg	[15:0]	RDATA;

initial
begin
   RDATA = $random;
end

// Look at the rising edge of the clock

always @ (posedge RCLK_g)
begin
	if	(RE)
	begin
		-> Read_e;
		if	(Time_Collision_Detected & Address_Collision_Detected) 
			RDATA <= 16'hXXXX;
		else
			for	(i=0;i<=BUS_WIDTH-1;i=i+1)
				RDATA[i]	<= Memory[RADDR*BUS_WIDTH+i];
	end
end

`ifdef TIMINGCHECK
specify
   (RCLK *> RDATA[0]) = (1.0, 1.0);
   (RCLK *> RDATA[1]) = (1.0, 1.0);
   (RCLK *> RDATA[2]) = (1.0, 1.0);
   (RCLK *> RDATA[3]) = (1.0, 1.0);
   (RCLK *> RDATA[4]) = (1.0, 1.0);
   (RCLK *> RDATA[5]) = (1.0, 1.0);
   (RCLK *> RDATA[6]) = (1.0, 1.0);
   (RCLK *> RDATA[7]) = (1.0, 1.0);
   (RCLK *> RDATA[8]) = (1.0, 1.0);
   (RCLK *> RDATA[9]) = (1.0, 1.0);
   (RCLK *> RDATA[10]) = (1.0, 1.0);
   (RCLK *> RDATA[11]) = (1.0, 1.0);
   (RCLK *> RDATA[12]) = (1.0, 1.0);
   (RCLK *> RDATA[13]) = (1.0, 1.0);
   (RCLK *> RDATA[14]) = (1.0, 1.0);
   (RCLK *> RDATA[15]) = (1.0, 1.0);
   $setup(posedge MASK[0], posedge WCLK, 1.0);
   $setup(negedge MASK[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[0], 1.0);
   $hold(posedge WCLK, negedge MASK[0], 1.0);
   $setup(posedge MASK[1], posedge WCLK, 1.0);
   $setup(negedge MASK[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[1], 1.0);
   $hold(posedge WCLK, negedge MASK[1], 1.0);
   $setup(posedge MASK[2], posedge WCLK, 1.0);
   $setup(negedge MASK[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[2], 1.0);
   $hold(posedge WCLK, negedge MASK[2], 1.0);
   $setup(posedge MASK[3], posedge WCLK, 1.0);
   $setup(negedge MASK[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[3], 1.0);
   $hold(posedge WCLK, negedge MASK[3], 1.0);
   $setup(posedge MASK[4], posedge WCLK, 1.0);
   $setup(negedge MASK[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[4], 1.0);
   $hold(posedge WCLK, negedge MASK[4], 1.0);
   $setup(posedge MASK[5], posedge WCLK, 1.0);
   $setup(negedge MASK[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[5], 1.0);
   $hold(posedge WCLK, negedge MASK[5], 1.0);
   $setup(posedge MASK[6], posedge WCLK, 1.0);
   $setup(negedge MASK[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[6], 1.0);
   $hold(posedge WCLK, negedge MASK[6], 1.0);
   $setup(posedge MASK[7], posedge WCLK, 1.0);
   $setup(negedge MASK[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[7], 1.0);
   $hold(posedge WCLK, negedge MASK[7], 1.0);
   $setup(posedge MASK[8], posedge WCLK, 1.0);
   $setup(negedge MASK[8], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[8], 1.0);
   $hold(posedge WCLK, negedge MASK[8], 1.0);
   $setup(posedge MASK[9], posedge WCLK, 1.0);
   $setup(negedge MASK[9], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[9], 1.0);
   $hold(posedge WCLK, negedge MASK[9], 1.0);
   $setup(posedge MASK[10], posedge WCLK, 1.0);
   $setup(negedge MASK[10], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[10], 1.0);
   $hold(posedge WCLK, negedge MASK[10], 1.0);
   $setup(posedge MASK[11], posedge WCLK, 1.0);
   $setup(negedge MASK[11], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[11], 1.0);
   $hold(posedge WCLK, negedge MASK[11], 1.0);
   $setup(posedge MASK[12], posedge WCLK, 1.0);
   $setup(negedge MASK[12], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[12], 1.0);
   $hold(posedge WCLK, negedge MASK[12], 1.0);
   $setup(posedge MASK[13], posedge WCLK, 1.0);
   $setup(negedge MASK[13], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[13], 1.0);
   $hold(posedge WCLK, negedge MASK[13], 1.0);
   $setup(posedge MASK[14], posedge WCLK, 1.0);
   $setup(negedge MASK[14], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[14], 1.0);
   $hold(posedge WCLK, negedge MASK[14], 1.0);
   $setup(posedge MASK[15], posedge WCLK, 1.0);
   $setup(negedge MASK[15], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[15], 1.0);
   $hold(posedge WCLK, negedge MASK[15], 1.0);
   $setup(posedge WADDR[0], posedge WCLK, 1.0);
   $setup(negedge WADDR[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[0], 1.0);
   $hold(posedge WCLK, negedge WADDR[0], 1.0);
   $setup(posedge WADDR[1], posedge WCLK, 1.0);
   $setup(negedge WADDR[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[1], 1.0);
   $hold(posedge WCLK, negedge WADDR[1], 1.0);
   $setup(posedge WADDR[2], posedge WCLK, 1.0);
   $setup(negedge WADDR[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[2], 1.0);
   $hold(posedge WCLK, negedge WADDR[2], 1.0);
   $setup(posedge WADDR[3], posedge WCLK, 1.0);
   $setup(negedge WADDR[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[3], 1.0);
   $hold(posedge WCLK, negedge WADDR[3], 1.0);
   $setup(posedge WADDR[4], posedge WCLK, 1.0);
   $setup(negedge WADDR[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[4], 1.0);
   $hold(posedge WCLK, negedge WADDR[4], 1.0);
   $setup(posedge WADDR[5], posedge WCLK, 1.0);
   $setup(negedge WADDR[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[5], 1.0);
   $hold(posedge WCLK, negedge WADDR[5], 1.0);
   $setup(posedge WADDR[6], posedge WCLK, 1.0);
   $setup(negedge WADDR[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[6], 1.0);
   $hold(posedge WCLK, negedge WADDR[6], 1.0);
   $setup(posedge WADDR[7], posedge WCLK, 1.0);
   $setup(negedge WADDR[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[7], 1.0);
   $hold(posedge WCLK, negedge WADDR[7], 1.0);
   $setup(posedge WDATA[0], posedge WCLK, 1.0);
   $setup(negedge WDATA[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[0], 1.0);
   $hold(posedge WCLK, negedge WDATA[0], 1.0);
   $setup(posedge WDATA[1], posedge WCLK, 1.0);
   $setup(negedge WDATA[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[1], 1.0);
   $hold(posedge WCLK, negedge WDATA[1], 1.0);
   $setup(posedge WDATA[2], posedge WCLK, 1.0);
   $setup(negedge WDATA[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[2], 1.0);
   $hold(posedge WCLK, negedge WDATA[2], 1.0);
   $setup(posedge WDATA[3], posedge WCLK, 1.0);
   $setup(negedge WDATA[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[3], 1.0);
   $hold(posedge WCLK, negedge WDATA[3], 1.0);
   $setup(posedge WDATA[4], posedge WCLK, 1.0);
   $setup(negedge WDATA[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[4], 1.0);
   $hold(posedge WCLK, negedge WDATA[4], 1.0);
   $setup(posedge WDATA[5], posedge WCLK, 1.0);
   $setup(negedge WDATA[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[5], 1.0);
   $hold(posedge WCLK, negedge WDATA[5], 1.0);
   $setup(posedge WDATA[6], posedge WCLK, 1.0);
   $setup(negedge WDATA[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[6], 1.0);
   $hold(posedge WCLK, negedge WDATA[6], 1.0);
   $setup(posedge WDATA[7], posedge WCLK, 1.0);
   $setup(negedge WDATA[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[7], 1.0);
   $hold(posedge WCLK, negedge WDATA[7], 1.0);
   $setup(posedge WDATA[8], posedge WCLK, 1.0);
   $setup(negedge WDATA[8], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[8], 1.0);
   $hold(posedge WCLK, negedge WDATA[8], 1.0);
   $setup(posedge WDATA[9], posedge WCLK, 1.0);
   $setup(negedge WDATA[9], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[9], 1.0);
   $hold(posedge WCLK, negedge WDATA[9], 1.0);
   $setup(posedge WDATA[10], posedge WCLK, 1.0);
   $setup(negedge WDATA[10], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[10], 1.0);
   $hold(posedge WCLK, negedge WDATA[10], 1.0);
   $setup(posedge WDATA[11], posedge WCLK, 1.0);
   $setup(negedge WDATA[11], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[11], 1.0);
   $hold(posedge WCLK, negedge WDATA[11], 1.0);
   $setup(posedge WDATA[12], posedge WCLK, 1.0);
   $setup(negedge WDATA[12], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[12], 1.0);
   $hold(posedge WCLK, negedge WDATA[12], 1.0);
   $setup(posedge WDATA[13], posedge WCLK, 1.0);
   $setup(negedge WDATA[13], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[13], 1.0);
   $hold(posedge WCLK, negedge WDATA[13], 1.0);
   $setup(posedge WDATA[14], posedge WCLK, 1.0);
   $setup(negedge WDATA[14], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[14], 1.0);
   $hold(posedge WCLK, negedge WDATA[14], 1.0);
   $setup(posedge WDATA[15], posedge WCLK, 1.0);
   $setup(negedge WDATA[15], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[15], 1.0);
   $hold(posedge WCLK, negedge WDATA[15], 1.0);
   $setup(posedge WCLKE, posedge WCLK, 1.0);
   $setup(negedge WCLKE, posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WCLKE, 1.0);
   $hold(posedge WCLK, negedge WCLKE, 1.0);
   $setup(posedge WE, posedge WCLK, 1.0);
   $setup(negedge WE, posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WE, 1.0);
   $hold(posedge WCLK, negedge WE, 1.0);
   $setup(posedge RADDR[0], posedge RCLK, 1.0);
   $setup(negedge RADDR[0], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[0], 1.0);
   $hold(posedge RCLK, negedge RADDR[0], 1.0);
   $setup(posedge RADDR[1], posedge RCLK, 1.0);
   $setup(negedge RADDR[1], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[1], 1.0);
   $hold(posedge RCLK, negedge RADDR[1], 1.0);
   $setup(posedge RADDR[2], posedge RCLK, 1.0);
   $setup(negedge RADDR[2], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[2], 1.0);
   $hold(posedge RCLK, negedge RADDR[2], 1.0);
   $setup(posedge RADDR[3], posedge RCLK, 1.0);
   $setup(negedge RADDR[3], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[3], 1.0);
   $hold(posedge RCLK, negedge RADDR[3], 1.0);
   $setup(posedge RADDR[4], posedge RCLK, 1.0);
   $setup(negedge RADDR[4], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[4], 1.0);
   $hold(posedge RCLK, negedge RADDR[4], 1.0);
   $setup(posedge RADDR[5], posedge RCLK, 1.0);
   $setup(negedge RADDR[5], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[5], 1.0);
   $hold(posedge RCLK, negedge RADDR[5], 1.0);
   $setup(posedge RADDR[6], posedge RCLK, 1.0);
   $setup(negedge RADDR[6], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[6], 1.0);
   $hold(posedge RCLK, negedge RADDR[6], 1.0);
   $setup(posedge RADDR[7], posedge RCLK, 1.0);
   $setup(negedge RADDR[7], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[7], 1.0);
   $hold(posedge RCLK, negedge RADDR[7], 1.0);
   $setup(posedge RCLKE, posedge RCLK, 1.0);
   $setup(negedge RCLKE, posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RCLKE, 1.0);
   $hold(posedge RCLK, negedge RCLKE, 1.0);
   $setup(posedge RE, posedge RCLK, 1.0);
   $setup(negedge RE, posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RE, 1.0);
   $hold(posedge RCLK, negedge RE, 1.0);

endspecify
`endif

endmodule //SB_RAM256x16

`timescale 1ps/1ps
module SB_RAM256x16NR (RDATA, RCLKN, RCLKE, RE, RADDR, WCLK, WCLKE, WE, WADDR, MASK, WDATA);
output [15:0] RDATA;
input RCLKN;
input RCLKE;
input RE;
input [7:0] RADDR;
input WCLK;
input WCLKE;
input WE;
input [7:0] WADDR;
input [15:0] MASK;
input [15:0] WDATA;

parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

wire RCLK;
assign (weak0, weak1) RCLKE =1'b1 ;
assign (weak0, weak1) RE =1'b0 ;
assign (weak0, weak1) WCLKE =1'b1 ;
assign (weak0, weak1) WE =1'b0 ;
assign RCLK = ~RCLKN;

SB_RAM256x16 sb_ram256X16r_inst (
	.RDATA(RDATA),
	.RCLK(RCLK),
	.RCLKE(RCLKE),
	.RE(RE),
	.RADDR(RADDR),
	.WCLK(WCLK),
	.WCLKE(WCLKE),
	.WE(WE),
	.WADDR(WADDR),
	.MASK(MASK),
	.WDATA(WDATA));

defparam sb_ram256X16r_inst.INIT_0 = INIT_0;
defparam sb_ram256X16r_inst.INIT_1 = INIT_1;
defparam sb_ram256X16r_inst.INIT_2 = INIT_2;
defparam sb_ram256X16r_inst.INIT_3 = INIT_3;
defparam sb_ram256X16r_inst.INIT_4 = INIT_4;
defparam sb_ram256X16r_inst.INIT_5 = INIT_5;
defparam sb_ram256X16r_inst.INIT_6 = INIT_6;
defparam sb_ram256X16r_inst.INIT_7 = INIT_7;
defparam sb_ram256X16r_inst.INIT_8 = INIT_8;
defparam sb_ram256X16r_inst.INIT_9 = INIT_9;
defparam sb_ram256X16r_inst.INIT_A = INIT_A;
defparam sb_ram256X16r_inst.INIT_B = INIT_B;
defparam sb_ram256X16r_inst.INIT_C = INIT_C;
defparam sb_ram256X16r_inst.INIT_D = INIT_D;
defparam sb_ram256X16r_inst.INIT_E = INIT_E;
defparam sb_ram256X16r_inst.INIT_F = INIT_F;

`ifdef TIMINGCHECK
specify
   (RCLKN *> RDATA[0]) = (1.0, 1.0);
   (RCLKN *> RDATA[1]) = (1.0, 1.0);
   (RCLKN *> RDATA[2]) = (1.0, 1.0);
   (RCLKN *> RDATA[3]) = (1.0, 1.0);
   (RCLKN *> RDATA[4]) = (1.0, 1.0);
   (RCLKN *> RDATA[5]) = (1.0, 1.0);
   (RCLKN *> RDATA[6]) = (1.0, 1.0);
   (RCLKN *> RDATA[7]) = (1.0, 1.0);
   (RCLKN *> RDATA[8]) = (1.0, 1.0);
   (RCLKN *> RDATA[9]) = (1.0, 1.0);
   (RCLKN *> RDATA[10]) = (1.0, 1.0);
   (RCLKN *> RDATA[11]) = (1.0, 1.0);
   (RCLKN *> RDATA[12]) = (1.0, 1.0);
   (RCLKN *> RDATA[13]) = (1.0, 1.0);
   (RCLKN *> RDATA[14]) = (1.0, 1.0);
   (RCLKN *> RDATA[15]) = (1.0, 1.0);
   $setup(posedge MASK[0], posedge WCLK, 1.0);
   $setup(negedge MASK[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[0], 1.0);
   $hold(posedge WCLK, negedge MASK[0], 1.0);
   $setup(posedge MASK[1], posedge WCLK, 1.0);
   $setup(negedge MASK[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[1], 1.0);
   $hold(posedge WCLK, negedge MASK[1], 1.0);
   $setup(posedge MASK[2], posedge WCLK, 1.0);
   $setup(negedge MASK[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[2], 1.0);
   $hold(posedge WCLK, negedge MASK[2], 1.0);
   $setup(posedge MASK[3], posedge WCLK, 1.0);
   $setup(negedge MASK[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[3], 1.0);
   $hold(posedge WCLK, negedge MASK[3], 1.0);
   $setup(posedge MASK[4], posedge WCLK, 1.0);
   $setup(negedge MASK[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[4], 1.0);
   $hold(posedge WCLK, negedge MASK[4], 1.0);
   $setup(posedge MASK[5], posedge WCLK, 1.0);
   $setup(negedge MASK[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[5], 1.0);
   $hold(posedge WCLK, negedge MASK[5], 1.0);
   $setup(posedge MASK[6], posedge WCLK, 1.0);
   $setup(negedge MASK[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[6], 1.0);
   $hold(posedge WCLK, negedge MASK[6], 1.0);
   $setup(posedge MASK[7], posedge WCLK, 1.0);
   $setup(negedge MASK[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[7], 1.0);
   $hold(posedge WCLK, negedge MASK[7], 1.0);
   $setup(posedge MASK[8], posedge WCLK, 1.0);
   $setup(negedge MASK[8], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[8], 1.0);
   $hold(posedge WCLK, negedge MASK[8], 1.0);
   $setup(posedge MASK[9], posedge WCLK, 1.0);
   $setup(negedge MASK[9], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[9], 1.0);
   $hold(posedge WCLK, negedge MASK[9], 1.0);
   $setup(posedge MASK[10], posedge WCLK, 1.0);
   $setup(negedge MASK[10], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[10], 1.0);
   $hold(posedge WCLK, negedge MASK[10], 1.0);
   $setup(posedge MASK[11], posedge WCLK, 1.0);
   $setup(negedge MASK[11], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[11], 1.0);
   $hold(posedge WCLK, negedge MASK[11], 1.0);
   $setup(posedge MASK[12], posedge WCLK, 1.0);
   $setup(negedge MASK[12], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[12], 1.0);
   $hold(posedge WCLK, negedge MASK[12], 1.0);
   $setup(posedge MASK[13], posedge WCLK, 1.0);
   $setup(negedge MASK[13], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[13], 1.0);
   $hold(posedge WCLK, negedge MASK[13], 1.0);
   $setup(posedge MASK[14], posedge WCLK, 1.0);
   $setup(negedge MASK[14], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[14], 1.0);
   $hold(posedge WCLK, negedge MASK[14], 1.0);
   $setup(posedge MASK[15], posedge WCLK, 1.0);
   $setup(negedge MASK[15], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[15], 1.0);
   $hold(posedge WCLK, negedge MASK[15], 1.0);
   $setup(posedge WADDR[0], posedge WCLK, 1.0);
   $setup(negedge WADDR[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[0], 1.0);
   $hold(posedge WCLK, negedge WADDR[0], 1.0);
   $setup(posedge WADDR[1], posedge WCLK, 1.0);
   $setup(negedge WADDR[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[1], 1.0);
   $hold(posedge WCLK, negedge WADDR[1], 1.0);
   $setup(posedge WADDR[2], posedge WCLK, 1.0);
   $setup(negedge WADDR[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[2], 1.0);
   $hold(posedge WCLK, negedge WADDR[2], 1.0);
   $setup(posedge WADDR[3], posedge WCLK, 1.0);
   $setup(negedge WADDR[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[3], 1.0);
   $hold(posedge WCLK, negedge WADDR[3], 1.0);
   $setup(posedge WADDR[4], posedge WCLK, 1.0);
   $setup(negedge WADDR[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[4], 1.0);
   $hold(posedge WCLK, negedge WADDR[4], 1.0);
   $setup(posedge WADDR[5], posedge WCLK, 1.0);
   $setup(negedge WADDR[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[5], 1.0);
   $hold(posedge WCLK, negedge WADDR[5], 1.0);
   $setup(posedge WADDR[6], posedge WCLK, 1.0);
   $setup(negedge WADDR[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[6], 1.0);
   $hold(posedge WCLK, negedge WADDR[6], 1.0);
   $setup(posedge WADDR[7], posedge WCLK, 1.0);
   $setup(negedge WADDR[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[7], 1.0);
   $hold(posedge WCLK, negedge WADDR[7], 1.0);
   $setup(posedge WDATA[0], posedge WCLK, 1.0);
   $setup(negedge WDATA[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[0], 1.0);
   $hold(posedge WCLK, negedge WDATA[0], 1.0);
   $setup(posedge WDATA[1], posedge WCLK, 1.0);
   $setup(negedge WDATA[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[1], 1.0);
   $hold(posedge WCLK, negedge WDATA[1], 1.0);
   $setup(posedge WDATA[2], posedge WCLK, 1.0);
   $setup(negedge WDATA[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[2], 1.0);
   $hold(posedge WCLK, negedge WDATA[2], 1.0);
   $setup(posedge WDATA[3], posedge WCLK, 1.0);
   $setup(negedge WDATA[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[3], 1.0);
   $hold(posedge WCLK, negedge WDATA[3], 1.0);
   $setup(posedge WDATA[4], posedge WCLK, 1.0);
   $setup(negedge WDATA[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[4], 1.0);
   $hold(posedge WCLK, negedge WDATA[4], 1.0);
   $setup(posedge WDATA[5], posedge WCLK, 1.0);
   $setup(negedge WDATA[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[5], 1.0);
   $hold(posedge WCLK, negedge WDATA[5], 1.0);
   $setup(posedge WDATA[6], posedge WCLK, 1.0);
   $setup(negedge WDATA[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[6], 1.0);
   $hold(posedge WCLK, negedge WDATA[6], 1.0);
   $setup(posedge WDATA[7], posedge WCLK, 1.0);
   $setup(negedge WDATA[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[7], 1.0);
   $hold(posedge WCLK, negedge WDATA[7], 1.0);
   $setup(posedge WDATA[8], posedge WCLK, 1.0);
   $setup(negedge WDATA[8], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[8], 1.0);
   $hold(posedge WCLK, negedge WDATA[8], 1.0);
   $setup(posedge WDATA[9], posedge WCLK, 1.0);
   $setup(negedge WDATA[9], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[9], 1.0);
   $hold(posedge WCLK, negedge WDATA[9], 1.0);
   $setup(posedge WDATA[10], posedge WCLK, 1.0);
   $setup(negedge WDATA[10], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[10], 1.0);
   $hold(posedge WCLK, negedge WDATA[10], 1.0);
   $setup(posedge WDATA[11], posedge WCLK, 1.0);
   $setup(negedge WDATA[11], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[11], 1.0);
   $hold(posedge WCLK, negedge WDATA[11], 1.0);
   $setup(posedge WDATA[12], posedge WCLK, 1.0);
   $setup(negedge WDATA[12], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[12], 1.0);
   $hold(posedge WCLK, negedge WDATA[12], 1.0);
   $setup(posedge WDATA[13], posedge WCLK, 1.0);
   $setup(negedge WDATA[13], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[13], 1.0);
   $hold(posedge WCLK, negedge WDATA[13], 1.0);
   $setup(posedge WDATA[14], posedge WCLK, 1.0);
   $setup(negedge WDATA[14], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[14], 1.0);
   $hold(posedge WCLK, negedge WDATA[14], 1.0);
   $setup(posedge WDATA[15], posedge WCLK, 1.0);
   $setup(negedge WDATA[15], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[15], 1.0);
   $hold(posedge WCLK, negedge WDATA[15], 1.0);
   $setup(posedge WCLKE, posedge WCLK, 1.0);
   $setup(negedge WCLKE, posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WCLKE, 1.0);
   $hold(posedge WCLK, negedge WCLKE, 1.0);
   $setup(posedge WE, posedge WCLK, 1.0);
   $setup(negedge WE, posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WE, 1.0);
   $hold(posedge WCLK, negedge WE, 1.0);
   $setup(posedge RADDR[0], posedge RCLKN, 1.0);
   $setup(negedge RADDR[0], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[0], 1.0);
   $hold(posedge RCLKN, negedge RADDR[0], 1.0);
   $setup(posedge RADDR[1], posedge RCLKN, 1.0);
   $setup(negedge RADDR[1], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[1], 1.0);
   $hold(posedge RCLKN, negedge RADDR[1], 1.0);
   $setup(posedge RADDR[2], posedge RCLKN, 1.0);
   $setup(negedge RADDR[2], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[2], 1.0);
   $hold(posedge RCLKN, negedge RADDR[2], 1.0);
   $setup(posedge RADDR[3], posedge RCLKN, 1.0);
   $setup(negedge RADDR[3], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[3], 1.0);
   $hold(posedge RCLKN, negedge RADDR[3], 1.0);
   $setup(posedge RADDR[4], posedge RCLKN, 1.0);
   $setup(negedge RADDR[4], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[4], 1.0);
   $hold(posedge RCLKN, negedge RADDR[4], 1.0);
   $setup(posedge RADDR[5], posedge RCLKN, 1.0);
   $setup(negedge RADDR[5], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[5], 1.0);
   $hold(posedge RCLKN, negedge RADDR[5], 1.0);
   $setup(posedge RADDR[6], posedge RCLKN, 1.0);
   $setup(negedge RADDR[6], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[6], 1.0);
   $hold(posedge RCLKN, negedge RADDR[6], 1.0);
   $setup(posedge RADDR[7], posedge RCLKN, 1.0);
   $setup(negedge RADDR[7], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[7], 1.0);
   $hold(posedge RCLKN, negedge RADDR[7], 1.0);
   $setup(posedge RCLKE, posedge RCLKN, 1.0);
   $setup(negedge RCLKE, posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RCLKE, 1.0);
   $hold(posedge RCLKN, negedge RCLKE, 1.0);
   $setup(posedge RE, posedge RCLKN, 1.0);
   $setup(negedge RE, posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RE, 1.0);
   $hold(posedge RCLKN, negedge RE, 1.0);
   $recovery(posedge RCLKN, posedge WCLK, 1.0);
   $recovery(negedge RCLKN, posedge WCLK, 1.0);
   $removal(posedge RCLKN, posedge WCLK, 1.0);
   $removal(negedge RCLKN, posedge WCLK, 1.0);
   $recovery(posedge WCLK, posedge RCLKN, 1.0);
   $recovery(negedge WCLK, posedge RCLKN, 1.0);
   $removal(posedge WCLK, posedge RCLKN, 1.0);
   $removal(negedge WCLK, posedge RCLKN, 1.0);

endspecify
`endif
endmodule //SB_RAM256x16NR

`timescale 1ps/1ps
module SB_RAM256x16NW (RDATA, RCLK, RCLKE, RE, RADDR, WCLKN, WCLKE, WE, WADDR, MASK, WDATA);
output [15:0] RDATA;
input RCLK;
input RCLKE;
input RE;
input [7:0] RADDR;
input WCLKN;
input WCLKE;
input WE;
input [7:0] WADDR;
input [15:0] MASK;
input [15:0] WDATA;

parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

wire WCLK;
assign (weak0, weak1) RCLKE =1'b1 ;
assign (weak0, weak1) RE =1'b0 ;
assign (weak0, weak1) WCLKE =1'b1 ;
assign (weak0, weak1) WE =1'b0 ;
assign WCLK = ~WCLKN;

SB_RAM256x16 sb_ram256X16w_inst (
	.RDATA(RDATA),
	.RCLK(RCLK),
	.RCLKE(RCLKE),
	.RE(RE),
	.RADDR(RADDR),
	.WCLK(WCLK),
	.WCLKE(WCLKE),
	.WE(WE),
	.WADDR(WADDR),
	.MASK(MASK),
	.WDATA(WDATA));

defparam sb_ram256X16w_inst.INIT_0 = INIT_0;
defparam sb_ram256X16w_inst.INIT_1 = INIT_1;
defparam sb_ram256X16w_inst.INIT_2 = INIT_2;
defparam sb_ram256X16w_inst.INIT_3 = INIT_3;
defparam sb_ram256X16w_inst.INIT_4 = INIT_4;
defparam sb_ram256X16w_inst.INIT_5 = INIT_5;
defparam sb_ram256X16w_inst.INIT_6 = INIT_6;
defparam sb_ram256X16w_inst.INIT_7 = INIT_7;
defparam sb_ram256X16w_inst.INIT_8 = INIT_8;
defparam sb_ram256X16w_inst.INIT_9 = INIT_9;
defparam sb_ram256X16w_inst.INIT_A = INIT_A;
defparam sb_ram256X16w_inst.INIT_B = INIT_B;
defparam sb_ram256X16w_inst.INIT_C = INIT_C;
defparam sb_ram256X16w_inst.INIT_D = INIT_D;
defparam sb_ram256X16w_inst.INIT_E = INIT_E;
defparam sb_ram256X16w_inst.INIT_F = INIT_F;

`ifdef TIMINGCHECK
specify
   (RCLK *> RDATA[0]) = (1.0, 1.0);
   (RCLK *> RDATA[1]) = (1.0, 1.0);
   (RCLK *> RDATA[2]) = (1.0, 1.0);
   (RCLK *> RDATA[3]) = (1.0, 1.0);
   (RCLK *> RDATA[4]) = (1.0, 1.0);
   (RCLK *> RDATA[5]) = (1.0, 1.0);
   (RCLK *> RDATA[6]) = (1.0, 1.0);
   (RCLK *> RDATA[7]) = (1.0, 1.0);
   (RCLK *> RDATA[8]) = (1.0, 1.0);
   (RCLK *> RDATA[9]) = (1.0, 1.0);
   (RCLK *> RDATA[10]) = (1.0, 1.0);
   (RCLK *> RDATA[11]) = (1.0, 1.0);
   (RCLK *> RDATA[12]) = (1.0, 1.0);
   (RCLK *> RDATA[13]) = (1.0, 1.0);
   (RCLK *> RDATA[14]) = (1.0, 1.0);
   (RCLK *> RDATA[15]) = (1.0, 1.0);
   $setup(posedge MASK[0], posedge WCLKN, 1.0);
   $setup(negedge MASK[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[0], 1.0);
   $hold(posedge WCLKN, negedge MASK[0], 1.0);
   $setup(posedge MASK[1], posedge WCLKN, 1.0);
   $setup(negedge MASK[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[1], 1.0);
   $hold(posedge WCLKN, negedge MASK[1], 1.0);
   $setup(posedge MASK[2], posedge WCLKN, 1.0);
   $setup(negedge MASK[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[2], 1.0);
   $hold(posedge WCLKN, negedge MASK[2], 1.0);
   $setup(posedge MASK[3], posedge WCLKN, 1.0);
   $setup(negedge MASK[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[3], 1.0);
   $hold(posedge WCLKN, negedge MASK[3], 1.0);
   $setup(posedge MASK[4], posedge WCLKN, 1.0);
   $setup(negedge MASK[4], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[4], 1.0);
   $hold(posedge WCLKN, negedge MASK[4], 1.0);
   $setup(posedge MASK[5], posedge WCLKN, 1.0);
   $setup(negedge MASK[5], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[5], 1.0);
   $hold(posedge WCLKN, negedge MASK[5], 1.0);
   $setup(posedge MASK[6], posedge WCLKN, 1.0);
   $setup(negedge MASK[6], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[6], 1.0);
   $hold(posedge WCLKN, negedge MASK[6], 1.0);
   $setup(posedge MASK[7], posedge WCLKN, 1.0);
   $setup(negedge MASK[7], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[7], 1.0);
   $hold(posedge WCLKN, negedge MASK[7], 1.0);
   $setup(posedge MASK[8], posedge WCLKN, 1.0);
   $setup(negedge MASK[8], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[8], 1.0);
   $hold(posedge WCLKN, negedge MASK[8], 1.0);
   $setup(posedge MASK[9], posedge WCLKN, 1.0);
   $setup(negedge MASK[9], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[9], 1.0);
   $hold(posedge WCLKN, negedge MASK[9], 1.0);
   $setup(posedge MASK[10], posedge WCLKN, 1.0);
   $setup(negedge MASK[10], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[10], 1.0);
   $hold(posedge WCLKN, negedge MASK[10], 1.0);
   $setup(posedge MASK[11], posedge WCLKN, 1.0);
   $setup(negedge MASK[11], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[11], 1.0);
   $hold(posedge WCLKN, negedge MASK[11], 1.0);
   $setup(posedge MASK[12], posedge WCLKN, 1.0);
   $setup(negedge MASK[12], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[12], 1.0);
   $hold(posedge WCLKN, negedge MASK[12], 1.0);
   $setup(posedge MASK[13], posedge WCLKN, 1.0);
   $setup(negedge MASK[13], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[13], 1.0);
   $hold(posedge WCLKN, negedge MASK[13], 1.0);
   $setup(posedge MASK[14], posedge WCLKN, 1.0);
   $setup(negedge MASK[14], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[14], 1.0);
   $hold(posedge WCLKN, negedge MASK[14], 1.0);
   $setup(posedge MASK[15], posedge WCLKN, 1.0);
   $setup(negedge MASK[15], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[15], 1.0);
   $hold(posedge WCLKN, negedge MASK[15], 1.0);
   $setup(posedge WADDR[0], posedge WCLKN, 1.0);
   $setup(negedge WADDR[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[0], 1.0);
   $hold(posedge WCLKN, negedge WADDR[0], 1.0);
   $setup(posedge WADDR[1], posedge WCLKN, 1.0);
   $setup(negedge WADDR[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[1], 1.0);
   $hold(posedge WCLKN, negedge WADDR[1], 1.0);
   $setup(posedge WADDR[2], posedge WCLKN, 1.0);
   $setup(negedge WADDR[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[2], 1.0);
   $hold(posedge WCLKN, negedge WADDR[2], 1.0);
   $setup(posedge WADDR[3], posedge WCLKN, 1.0);
   $setup(negedge WADDR[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[3], 1.0);
   $hold(posedge WCLKN, negedge WADDR[3], 1.0);
   $setup(posedge WADDR[4], posedge WCLKN, 1.0);
   $setup(negedge WADDR[4], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[4], 1.0);
   $hold(posedge WCLKN, negedge WADDR[4], 1.0);
   $setup(posedge WADDR[5], posedge WCLKN, 1.0);
   $setup(negedge WADDR[5], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[5], 1.0);
   $hold(posedge WCLKN, negedge WADDR[5], 1.0);
   $setup(posedge WADDR[6], posedge WCLKN, 1.0);
   $setup(negedge WADDR[6], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[6], 1.0);
   $hold(posedge WCLKN, negedge WADDR[6], 1.0);
   $setup(posedge WADDR[7], posedge WCLKN, 1.0);
   $setup(negedge WADDR[7], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[7], 1.0);
   $hold(posedge WCLKN, negedge WADDR[7], 1.0);
   $setup(posedge WDATA[0], posedge WCLKN, 1.0);
   $setup(negedge WDATA[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[0], 1.0);
   $hold(posedge WCLKN, negedge WDATA[0], 1.0);
   $setup(posedge WDATA[1], posedge WCLKN, 1.0);
   $setup(negedge WDATA[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[1], 1.0);
   $hold(posedge WCLKN, negedge WDATA[1], 1.0);
   $setup(posedge WDATA[2], posedge WCLKN, 1.0);
   $setup(negedge WDATA[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[2], 1.0);
   $hold(posedge WCLKN, negedge WDATA[2], 1.0);
   $setup(posedge WDATA[3], posedge WCLKN, 1.0);
   $setup(negedge WDATA[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[3], 1.0);
   $hold(posedge WCLKN, negedge WDATA[3], 1.0);
   $setup(posedge WDATA[4], posedge WCLKN, 1.0);
   $setup(negedge WDATA[4], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[4], 1.0);
   $hold(posedge WCLKN, negedge WDATA[4], 1.0);
   $setup(posedge WDATA[5], posedge WCLKN, 1.0);
   $setup(negedge WDATA[5], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[5], 1.0);
   $hold(posedge WCLKN, negedge WDATA[5], 1.0);
   $setup(posedge WDATA[6], posedge WCLKN, 1.0);
   $setup(negedge WDATA[6], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[6], 1.0);
   $hold(posedge WCLKN, negedge WDATA[6], 1.0);
   $setup(posedge WDATA[7], posedge WCLKN, 1.0);
   $setup(negedge WDATA[7], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[7], 1.0);
   $hold(posedge WCLKN, negedge WDATA[7], 1.0);
   $setup(posedge WDATA[8], posedge WCLKN, 1.0);
   $setup(negedge WDATA[8], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[8], 1.0);
   $hold(posedge WCLKN, negedge WDATA[8], 1.0);
   $setup(posedge WDATA[9], posedge WCLKN, 1.0);
   $setup(negedge WDATA[9], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[9], 1.0);
   $hold(posedge WCLKN, negedge WDATA[9], 1.0);
   $setup(posedge WDATA[10], posedge WCLKN, 1.0);
   $setup(negedge WDATA[10], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[10], 1.0);
   $hold(posedge WCLKN, negedge WDATA[10], 1.0);
   $setup(posedge WDATA[11], posedge WCLKN, 1.0);
   $setup(negedge WDATA[11], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[11], 1.0);
   $hold(posedge WCLKN, negedge WDATA[11], 1.0);
   $setup(posedge WDATA[12], posedge WCLKN, 1.0);
   $setup(negedge WDATA[12], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[12], 1.0);
   $hold(posedge WCLKN, negedge WDATA[12], 1.0);
   $setup(posedge WDATA[13], posedge WCLKN, 1.0);
   $setup(negedge WDATA[13], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[13], 1.0);
   $hold(posedge WCLKN, negedge WDATA[13], 1.0);
   $setup(posedge WDATA[14], posedge WCLKN, 1.0);
   $setup(negedge WDATA[14], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[14], 1.0);
   $hold(posedge WCLKN, negedge WDATA[14], 1.0);
   $setup(posedge WDATA[15], posedge WCLKN, 1.0);
   $setup(negedge WDATA[15], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[15], 1.0);
   $hold(posedge WCLKN, negedge WDATA[15], 1.0);
   $setup(posedge WCLKE, posedge WCLKN, 1.0);
   $setup(negedge WCLKE, posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WCLKE, 1.0);
   $hold(posedge WCLKN, negedge WCLKE, 1.0);
   $setup(posedge WE, posedge WCLKN, 1.0);
   $setup(negedge WE, posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WE, 1.0);
   $hold(posedge WCLKN, negedge WE, 1.0);
   $setup(posedge RADDR[0], posedge RCLK, 1.0);
   $setup(negedge RADDR[0], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[0], 1.0);
   $hold(posedge RCLK, negedge RADDR[0], 1.0);
   $setup(posedge RADDR[1], posedge RCLK, 1.0);
   $setup(negedge RADDR[1], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[1], 1.0);
   $hold(posedge RCLK, negedge RADDR[1], 1.0);
   $setup(posedge RADDR[2], posedge RCLK, 1.0);
   $setup(negedge RADDR[2], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[2], 1.0);
   $hold(posedge RCLK, negedge RADDR[2], 1.0);
   $setup(posedge RADDR[3], posedge RCLK, 1.0);
   $setup(negedge RADDR[3], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[3], 1.0);
   $hold(posedge RCLK, negedge RADDR[3], 1.0);
   $setup(posedge RADDR[4], posedge RCLK, 1.0);
   $setup(negedge RADDR[4], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[4], 1.0);
   $hold(posedge RCLK, negedge RADDR[4], 1.0);
   $setup(posedge RADDR[5], posedge RCLK, 1.0);
   $setup(negedge RADDR[5], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[5], 1.0);
   $hold(posedge RCLK, negedge RADDR[5], 1.0);
   $setup(posedge RADDR[6], posedge RCLK, 1.0);
   $setup(negedge RADDR[6], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[6], 1.0);
   $hold(posedge RCLK, negedge RADDR[6], 1.0);
   $setup(posedge RADDR[7], posedge RCLK, 1.0);
   $setup(negedge RADDR[7], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[7], 1.0);
   $hold(posedge RCLK, negedge RADDR[7], 1.0);
   $setup(posedge RCLKE, posedge RCLK, 1.0);
   $setup(negedge RCLKE, posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RCLKE, 1.0);
   $hold(posedge RCLK, negedge RCLKE, 1.0);
   $setup(posedge RE, posedge RCLK, 1.0);
   $setup(negedge RE, posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RE, 1.0);
   $hold(posedge RCLK, negedge RE, 1.0);
   $recovery(posedge RCLK, posedge WCLKN, 1.0);
   $recovery(negedge RCLK, posedge WCLKN, 1.0);
   $removal(posedge RCLK, posedge WCLKN, 1.0);
   $removal(negedge RCLK, posedge WCLKN, 1.0);
   $recovery(posedge WCLKN, posedge RCLK, 1.0);
   $recovery(negedge WCLKN, posedge RCLK, 1.0);
   $removal(posedge WCLKN, posedge RCLK, 1.0);
   $removal(negedge WCLKN, posedge RCLK, 1.0);

endspecify
`endif
endmodule //SB_RAM256x16NW

`timescale 1ps/1ps

module SB_RAM256x16NRNW (RDATA, RCLKN, RCLKE, RE, RADDR, WCLKN, WCLKE, WE, WADDR, MASK, WDATA);
output [15:0] RDATA;
input RCLKN;
input RCLKE;
input RE;
input [7:0] RADDR;
input WCLKN;
input WCLKE;
input WE;
input [7:0] WADDR;
input [15:0] MASK;
input [15:0] WDATA;

parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

wire RCLK, WCLK;
assign (weak0, weak1) RCLKE =1'b1 ;
assign (weak0, weak1) RE =1'b0 ;
assign (weak0, weak1) WCLKE =1'b1 ;
assign (weak0, weak1) WE =1'b0 ;
assign RCLK = ~RCLKN;
assign WCLK = ~WCLKN;

SB_RAM256x16 sb_ram256X16rw_inst (
	.RDATA(RDATA),
	.RCLK(RCLK),
	.RCLKE(RCLKE),
	.RE(RE),
	.RADDR(RADDR),
	.WCLK(WCLK),
	.WCLKE(WCLKE),
	.WE(WE),
	.WADDR(WADDR),
	.MASK(MASK),
	.WDATA(WDATA));

defparam sb_ram256X16rw_inst.INIT_0 = INIT_0;
defparam sb_ram256X16rw_inst.INIT_1 = INIT_1;
defparam sb_ram256X16rw_inst.INIT_2 = INIT_2;
defparam sb_ram256X16rw_inst.INIT_3 = INIT_3;
defparam sb_ram256X16rw_inst.INIT_4 = INIT_4;
defparam sb_ram256X16rw_inst.INIT_5 = INIT_5;
defparam sb_ram256X16rw_inst.INIT_6 = INIT_6;
defparam sb_ram256X16rw_inst.INIT_7 = INIT_7;
defparam sb_ram256X16rw_inst.INIT_8 = INIT_8;
defparam sb_ram256X16rw_inst.INIT_9 = INIT_9;
defparam sb_ram256X16rw_inst.INIT_A = INIT_A;
defparam sb_ram256X16rw_inst.INIT_B = INIT_B;
defparam sb_ram256X16rw_inst.INIT_C = INIT_C;
defparam sb_ram256X16rw_inst.INIT_D = INIT_D;
defparam sb_ram256X16rw_inst.INIT_E = INIT_E;
defparam sb_ram256X16rw_inst.INIT_F = INIT_F;

`ifdef TIMINGCHECK
specify
   (RCLKN *> RDATA[0]) = (1.0, 1.0);
   (RCLKN *> RDATA[1]) = (1.0, 1.0);
   (RCLKN *> RDATA[2]) = (1.0, 1.0);
   (RCLKN *> RDATA[3]) = (1.0, 1.0);
   (RCLKN *> RDATA[4]) = (1.0, 1.0);
   (RCLKN *> RDATA[5]) = (1.0, 1.0);
   (RCLKN *> RDATA[6]) = (1.0, 1.0);
   (RCLKN *> RDATA[7]) = (1.0, 1.0);
   (RCLKN *> RDATA[8]) = (1.0, 1.0);
   (RCLKN *> RDATA[9]) = (1.0, 1.0);
   (RCLKN *> RDATA[10]) = (1.0, 1.0);
   (RCLKN *> RDATA[11]) = (1.0, 1.0);
   (RCLKN *> RDATA[12]) = (1.0, 1.0);
   (RCLKN *> RDATA[13]) = (1.0, 1.0);
   (RCLKN *> RDATA[14]) = (1.0, 1.0);
   (RCLKN *> RDATA[15]) = (1.0, 1.0);
   $setup(posedge MASK[0], posedge WCLKN, 1.0);
   $setup(negedge MASK[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[0], 1.0);
   $hold(posedge WCLKN, negedge MASK[0], 1.0);
   $setup(posedge MASK[1], posedge WCLKN, 1.0);
   $setup(negedge MASK[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[1], 1.0);
   $hold(posedge WCLKN, negedge MASK[1], 1.0);
   $setup(posedge MASK[2], posedge WCLKN, 1.0);
   $setup(negedge MASK[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[2], 1.0);
   $hold(posedge WCLKN, negedge MASK[2], 1.0);
   $setup(posedge MASK[3], posedge WCLKN, 1.0);
   $setup(negedge MASK[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[3], 1.0);
   $hold(posedge WCLKN, negedge MASK[3], 1.0);
   $setup(posedge MASK[4], posedge WCLKN, 1.0);
   $setup(negedge MASK[4], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[4], 1.0);
   $hold(posedge WCLKN, negedge MASK[4], 1.0);
   $setup(posedge MASK[5], posedge WCLKN, 1.0);
   $setup(negedge MASK[5], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[5], 1.0);
   $hold(posedge WCLKN, negedge MASK[5], 1.0);
   $setup(posedge MASK[6], posedge WCLKN, 1.0);
   $setup(negedge MASK[6], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[6], 1.0);
   $hold(posedge WCLKN, negedge MASK[6], 1.0);
   $setup(posedge MASK[7], posedge WCLKN, 1.0);
   $setup(negedge MASK[7], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[7], 1.0);
   $hold(posedge WCLKN, negedge MASK[7], 1.0);
   $setup(posedge MASK[8], posedge WCLKN, 1.0);
   $setup(negedge MASK[8], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[8], 1.0);
   $hold(posedge WCLKN, negedge MASK[8], 1.0);
   $setup(posedge MASK[9], posedge WCLKN, 1.0);
   $setup(negedge MASK[9], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[9], 1.0);
   $hold(posedge WCLKN, negedge MASK[9], 1.0);
   $setup(posedge MASK[10], posedge WCLKN, 1.0);
   $setup(negedge MASK[10], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[10], 1.0);
   $hold(posedge WCLKN, negedge MASK[10], 1.0);
   $setup(posedge MASK[11], posedge WCLKN, 1.0);
   $setup(negedge MASK[11], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[11], 1.0);
   $hold(posedge WCLKN, negedge MASK[11], 1.0);
   $setup(posedge MASK[12], posedge WCLKN, 1.0);
   $setup(negedge MASK[12], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[12], 1.0);
   $hold(posedge WCLKN, negedge MASK[12], 1.0);
   $setup(posedge MASK[13], posedge WCLKN, 1.0);
   $setup(negedge MASK[13], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[13], 1.0);
   $hold(posedge WCLKN, negedge MASK[13], 1.0);
   $setup(posedge MASK[14], posedge WCLKN, 1.0);
   $setup(negedge MASK[14], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[14], 1.0);
   $hold(posedge WCLKN, negedge MASK[14], 1.0);
   $setup(posedge MASK[15], posedge WCLKN, 1.0);
   $setup(negedge MASK[15], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[15], 1.0);
   $hold(posedge WCLKN, negedge MASK[15], 1.0);
   $setup(posedge WADDR[0], posedge WCLKN, 1.0);
   $setup(negedge WADDR[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[0], 1.0);
   $hold(posedge WCLKN, negedge WADDR[0], 1.0);
   $setup(posedge WADDR[1], posedge WCLKN, 1.0);
   $setup(negedge WADDR[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[1], 1.0);
   $hold(posedge WCLKN, negedge WADDR[1], 1.0);
   $setup(posedge WADDR[2], posedge WCLKN, 1.0);
   $setup(negedge WADDR[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[2], 1.0);
   $hold(posedge WCLKN, negedge WADDR[2], 1.0);
   $setup(posedge WADDR[3], posedge WCLKN, 1.0);
   $setup(negedge WADDR[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[3], 1.0);
   $hold(posedge WCLKN, negedge WADDR[3], 1.0);
   $setup(posedge WADDR[4], posedge WCLKN, 1.0);
   $setup(negedge WADDR[4], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[4], 1.0);
   $hold(posedge WCLKN, negedge WADDR[4], 1.0);
   $setup(posedge WADDR[5], posedge WCLKN, 1.0);
   $setup(negedge WADDR[5], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[5], 1.0);
   $hold(posedge WCLKN, negedge WADDR[5], 1.0);
   $setup(posedge WADDR[6], posedge WCLKN, 1.0);
   $setup(negedge WADDR[6], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[6], 1.0);
   $hold(posedge WCLKN, negedge WADDR[6], 1.0);
   $setup(posedge WADDR[7], posedge WCLKN, 1.0);
   $setup(negedge WADDR[7], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[7], 1.0);
   $hold(posedge WCLKN, negedge WADDR[7], 1.0);
   $setup(posedge WDATA[0], posedge WCLKN, 1.0);
   $setup(negedge WDATA[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[0], 1.0);
   $hold(posedge WCLKN, negedge WDATA[0], 1.0);
   $setup(posedge WDATA[1], posedge WCLKN, 1.0);
   $setup(negedge WDATA[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[1], 1.0);
   $hold(posedge WCLKN, negedge WDATA[1], 1.0);
   $setup(posedge WDATA[2], posedge WCLKN, 1.0);
   $setup(negedge WDATA[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[2], 1.0);
   $hold(posedge WCLKN, negedge WDATA[2], 1.0);
   $setup(posedge WDATA[3], posedge WCLKN, 1.0);
   $setup(negedge WDATA[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[3], 1.0);
   $hold(posedge WCLKN, negedge WDATA[3], 1.0);
   $setup(posedge WDATA[4], posedge WCLKN, 1.0);
   $setup(negedge WDATA[4], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[4], 1.0);
   $hold(posedge WCLKN, negedge WDATA[4], 1.0);
   $setup(posedge WDATA[5], posedge WCLKN, 1.0);
   $setup(negedge WDATA[5], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[5], 1.0);
   $hold(posedge WCLKN, negedge WDATA[5], 1.0);
   $setup(posedge WDATA[6], posedge WCLKN, 1.0);
   $setup(negedge WDATA[6], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[6], 1.0);
   $hold(posedge WCLKN, negedge WDATA[6], 1.0);
   $setup(posedge WDATA[7], posedge WCLKN, 1.0);
   $setup(negedge WDATA[7], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[7], 1.0);
   $hold(posedge WCLKN, negedge WDATA[7], 1.0);
   $setup(posedge WDATA[8], posedge WCLKN, 1.0);
   $setup(negedge WDATA[8], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[8], 1.0);
   $hold(posedge WCLKN, negedge WDATA[8], 1.0);
   $setup(posedge WDATA[9], posedge WCLKN, 1.0);
   $setup(negedge WDATA[9], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[9], 1.0);
   $hold(posedge WCLKN, negedge WDATA[9], 1.0);
   $setup(posedge WDATA[10], posedge WCLKN, 1.0);
   $setup(negedge WDATA[10], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[10], 1.0);
   $hold(posedge WCLKN, negedge WDATA[10], 1.0);
   $setup(posedge WDATA[11], posedge WCLKN, 1.0);
   $setup(negedge WDATA[11], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[11], 1.0);
   $hold(posedge WCLKN, negedge WDATA[11], 1.0);
   $setup(posedge WDATA[12], posedge WCLKN, 1.0);
   $setup(negedge WDATA[12], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[12], 1.0);
   $hold(posedge WCLKN, negedge WDATA[12], 1.0);
   $setup(posedge WDATA[13], posedge WCLKN, 1.0);
   $setup(negedge WDATA[13], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[13], 1.0);
   $hold(posedge WCLKN, negedge WDATA[13], 1.0);
   $setup(posedge WDATA[14], posedge WCLKN, 1.0);
   $setup(negedge WDATA[14], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[14], 1.0);
   $hold(posedge WCLKN, negedge WDATA[14], 1.0);
   $setup(posedge WDATA[15], posedge WCLKN, 1.0);
   $setup(negedge WDATA[15], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[15], 1.0);
   $hold(posedge WCLKN, negedge WDATA[15], 1.0);
   $setup(posedge WCLKE, posedge WCLKN, 1.0);
   $setup(negedge WCLKE, posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WCLKE, 1.0);
   $hold(posedge WCLKN, negedge WCLKE, 1.0);
   $setup(posedge WE, posedge WCLKN, 1.0);
   $setup(negedge WE, posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WE, 1.0);
   $hold(posedge WCLKN, negedge WE, 1.0);
   $setup(posedge RADDR[0], posedge RCLKN, 1.0);
   $setup(negedge RADDR[0], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[0], 1.0);
   $hold(posedge RCLKN, negedge RADDR[0], 1.0);
   $setup(posedge RADDR[1], posedge RCLKN, 1.0);
   $setup(negedge RADDR[1], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[1], 1.0);
   $hold(posedge RCLKN, negedge RADDR[1], 1.0);
   $setup(posedge RADDR[2], posedge RCLKN, 1.0);
   $setup(negedge RADDR[2], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[2], 1.0);
   $hold(posedge RCLKN, negedge RADDR[2], 1.0);
   $setup(posedge RADDR[3], posedge RCLKN, 1.0);
   $setup(negedge RADDR[3], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[3], 1.0);
   $hold(posedge RCLKN, negedge RADDR[3], 1.0);
   $setup(posedge RADDR[4], posedge RCLKN, 1.0);
   $setup(negedge RADDR[4], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[4], 1.0);
   $hold(posedge RCLKN, negedge RADDR[4], 1.0);
   $setup(posedge RADDR[5], posedge RCLKN, 1.0);
   $setup(negedge RADDR[5], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[5], 1.0);
   $hold(posedge RCLKN, negedge RADDR[5], 1.0);
   $setup(posedge RADDR[6], posedge RCLKN, 1.0);
   $setup(negedge RADDR[6], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[6], 1.0);
   $hold(posedge RCLKN, negedge RADDR[6], 1.0);
   $setup(posedge RADDR[7], posedge RCLKN, 1.0);
   $setup(negedge RADDR[7], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[7], 1.0);
   $hold(posedge RCLKN, negedge RADDR[7], 1.0);
   $setup(posedge RCLKE, posedge RCLKN, 1.0);
   $setup(negedge RCLKE, posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RCLKE, 1.0);
   $hold(posedge RCLKN, negedge RCLKE, 1.0);
   $setup(posedge RE, posedge RCLKN, 1.0);
   $setup(negedge RE, posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RE, 1.0);
   $hold(posedge RCLKN, negedge RE, 1.0);
   $recovery(posedge RCLKN, posedge WCLKN, 1.0);
   $recovery(negedge RCLKN, posedge WCLKN, 1.0);
   $removal(posedge RCLKN, posedge WCLKN, 1.0);
   $removal(negedge RCLKN, posedge WCLKN, 1.0);
   $recovery(posedge WCLKN, posedge RCLKN, 1.0);
   $recovery(negedge WCLKN, posedge RCLKN, 1.0);
   $removal(posedge WCLKN, posedge RCLKN, 1.0);
   $removal(negedge WCLKN, posedge RCLKN, 1.0);

endspecify
`endif
endmodule //SB_RAM256x16NRNW

`timescale 1ps/1ps
module SB_RAM512x8 (RDATA, RCLK, RCLKE, RE, RADDR, WCLK, WCLKE, WE, WADDR, WDATA);
output [7:0] RDATA;
input RCLK;
input RCLKE;
input RE;
input [8:0] RADDR;
input WCLK;
input WCLKE;
input WE;
input [8:0] WADDR;
input [7:0] WDATA;

parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

// local Parameters
localparam			CLOCK_PERIOD = 200;	//
localparam 			DELAY	= (CLOCK_PERIOD/10);		// Clock-to-output delay. Zero
							// time delays can be confusing
							// and sometimes cause problems.
localparam 			BUS_WIDTH = 8;		// Width of RAM (number of bits)

localparam 			ADDRESS_BUS_SIZE = 9;	// Number of bits required to
							// represent the RAM address

localparam   ADDRESSABLE_SPACE  = 2**ADDRESS_BUS_SIZE;	// Decimal address range [2^Size:0]


// SIGNAL DECLARATIONS
wire			   	WCLK_g, RCLK_g;
reg 				WCLKE_sync, RCLKE_sync; 
assign (weak0, weak1) RCLKE =1'b1 ;
assign (weak0, weak1) RE =1'b0 ;
assign (weak0, weak1) WCLKE =1'b1 ;
assign (weak0, weak1) WE =1'b0 ;
reg	Memory	[BUS_WIDTH*ADDRESSABLE_SPACE-1:0];
// 
event Read_e, Write_e;

//////////////////// Collision detect begins here ///////////////////////////////
localparam 	TRUE = 1'b1;
localparam	FALSE = 1'b0;
reg 		Time_Collision_Detected = 1'b0;
wire		Address_Collision_Detected;

event Collision_e;

time COLLISION_TIME_WINDOW = (CLOCK_PERIOD/8); // This is an arbitray value, but is better than using an absolute 
						    // value, because the actual time window depends on the actual silicon 
						    // implementation. Thus the test is indicative of an Error and not
						    // guaranteed to be an error. Even so this is usefull.
time time_WCLK_RCLK, time_WCLK, time_RCLK;


//function reg Check_Timed_Window_Violation;
function	Check_Timed_Window_Violation;	//	by Jeffrey
input T1, T2, Minimum_Time_Window;
time T1, T2;
time Minimum_Time_Window;
time Difference;	
	begin
		Difference = (T1 - T2);
		if (Difference < 0) Difference = -Difference;
		Check_Timed_Window_Violation = (Difference < Minimum_Time_Window);
	end
endfunction


initial begin
       time_WCLK = CLOCK_PERIOD;	// Arbitrary initialisation value, ensure no window collison error on first clock edge.
       time_RCLK = (CLOCK_PERIOD*8);	// Arbitrary initialisation difference value, ensure no collision error on first clock edge.					
end

integer	i,j;


initial	//	initialize ram_4k by parameter, section by section
begin
	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[BUS_WIDTH*i+j]	=	INIT_0[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*1+BUS_WIDTH*i+j]	=	INIT_1[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*2+BUS_WIDTH*i+j]	=	INIT_2[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*3+BUS_WIDTH*i+j]	=	INIT_3[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*4+BUS_WIDTH*i+j]	=	INIT_4[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*5+BUS_WIDTH*i+j]	=	INIT_5[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*6+BUS_WIDTH*i+j]	=	INIT_6[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*7+BUS_WIDTH*i+j]	=	INIT_7[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*8+BUS_WIDTH*i+j]	=	INIT_8[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*9+BUS_WIDTH*i+j]	=	INIT_9[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*10+BUS_WIDTH*i+j]	=	INIT_A[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*11+BUS_WIDTH*i+j]	=	INIT_B[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*12+BUS_WIDTH*i+j]	=	INIT_C[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*13+BUS_WIDTH*i+j]	=	INIT_D[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*14+BUS_WIDTH*i+j]	=	INIT_E[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*15+BUS_WIDTH*i+j]	=	INIT_F[BUS_WIDTH*i+j];
	end

end

assign Address_Collision_Detected = ((RE & WE & WCLKE & RCLKE)&(WADDR == RADDR));


always @(WCLK or WCLKE) 
begin 
	if(~WCLK)
	WCLKE_sync = WCLKE;   	
end 

always @(RCLK or RCLKE) 
begin 
	if (~RCLK)
	RCLKE_sync = RCLKE; 	
end 

assign WCLK_g = WCLK & WCLKE_sync;
assign RCLK_g = RCLK & RCLKE_sync;
 
always @(posedge WCLK_g) begin
	time_WCLK = $time;
end

always @(posedge RCLK_g) begin
    	time_RCLK = $time;
end
integer	SB_RAM512X8_RDATA_log_file;					//.....................
initial	SB_RAM512X8_RDATA_log_file=("SB_RAM512X8_RDATA_log_file.txt");	//.....................
always @(posedge WCLK_g) begin

	Time_Collision_Detected = Check_Timed_Window_Violation(time_WCLK,time_RCLK,COLLISION_TIME_WINDOW);
        if (Time_Collision_Detected & Address_Collision_Detected)begin
        	$display("Warning: Write-Read collision detected, Data read value is XX\n");
 		$display("WCLK Time: %.3f   RCLK Time:%.3f  ",time_WCLK, time_RCLK,"WADDR: %d   RADDR:%d\n",WADDR, RADDR); 
 		$fdisplay(SB_RAM512X8_RDATA_log_file,"Warning: Write-Read collision detected, Data read value is XX\n");
		$fdisplay(SB_RAM512X8_RDATA_log_file,"WCLK Time: %.3f   RCLK Time:%.3f  ",time_WCLK, time_RCLK, "WADDR: %d   RADDR:%d\n",WADDR, RADDR); 	
 		-> Collision_e;
	end
end




//	code modify for universal verilog compiler

always @ (posedge WCLK_g)
begin
	if	(WE)
	begin
		-> Write_e;
		for	(i=0;i<=BUS_WIDTH-1; i=i+1)
		begin
			Memory[WADDR*BUS_WIDTH+i]	<=	WDATA[i];
		end
	end
end

//reg	[7:0]	RDATA = 0;
reg	[7:0]	RDATA;

initial
begin
   RDATA = $random;
end

// Look at the rising edge of the clock

always @ (posedge RCLK_g)
begin
	if	(RE)
	begin
		-> Read_e;
		if	(Time_Collision_Detected & Address_Collision_Detected) 
			RDATA <= 8'hXX;
		else
			for	(i=0;i<=BUS_WIDTH-1;i=i+1)
				RDATA[i]	<= Memory[RADDR*BUS_WIDTH+i];
	end
end

`ifdef TIMINGCHECK
specify
   (RCLK *> RDATA[0]) = (1.0, 1.0);
   (RCLK *> RDATA[1]) = (1.0, 1.0);
   (RCLK *> RDATA[2]) = (1.0, 1.0);
   (RCLK *> RDATA[3]) = (1.0, 1.0);
   (RCLK *> RDATA[4]) = (1.0, 1.0);
   (RCLK *> RDATA[5]) = (1.0, 1.0);
   (RCLK *> RDATA[6]) = (1.0, 1.0);
   (RCLK *> RDATA[7]) = (1.0, 1.0);
   $setup(posedge WADDR[0], posedge WCLK, 1.0);
   $setup(negedge WADDR[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[0], 1.0);
   $hold(posedge WCLK, negedge WADDR[0], 1.0);
   $setup(posedge WADDR[1], posedge WCLK, 1.0);
   $setup(negedge WADDR[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[1], 1.0);
   $hold(posedge WCLK, negedge WADDR[1], 1.0);
   $setup(posedge WADDR[2], posedge WCLK, 1.0);
   $setup(negedge WADDR[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[2], 1.0);
   $hold(posedge WCLK, negedge WADDR[2], 1.0);
   $setup(posedge WADDR[3], posedge WCLK, 1.0);
   $setup(negedge WADDR[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[3], 1.0);
   $hold(posedge WCLK, negedge WADDR[3], 1.0);
   $setup(posedge WADDR[4], posedge WCLK, 1.0);
   $setup(negedge WADDR[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[4], 1.0);
   $hold(posedge WCLK, negedge WADDR[4], 1.0);
   $setup(posedge WADDR[5], posedge WCLK, 1.0);
   $setup(negedge WADDR[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[5], 1.0);
   $hold(posedge WCLK, negedge WADDR[5], 1.0);
   $setup(posedge WADDR[6], posedge WCLK, 1.0);
   $setup(negedge WADDR[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[6], 1.0);
   $hold(posedge WCLK, negedge WADDR[6], 1.0);
   $setup(posedge WADDR[7], posedge WCLK, 1.0);
   $setup(negedge WADDR[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[7], 1.0);
   $hold(posedge WCLK, negedge WADDR[7], 1.0);
   $setup(posedge WADDR[8], posedge WCLK, 1.0);
   $setup(negedge WADDR[8], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[8], 1.0);
   $hold(posedge WCLK, negedge WADDR[8], 1.0);
   $setup(posedge WDATA[0], posedge WCLK, 1.0);
   $setup(negedge WDATA[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[0], 1.0);
   $hold(posedge WCLK, negedge WDATA[0], 1.0);
   $setup(posedge WDATA[1], posedge WCLK, 1.0);
   $setup(negedge WDATA[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[1], 1.0);
   $hold(posedge WCLK, negedge WDATA[1], 1.0);
   $setup(posedge WDATA[2], posedge WCLK, 1.0);
   $setup(negedge WDATA[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[2], 1.0);
   $hold(posedge WCLK, negedge WDATA[2], 1.0);
   $setup(posedge WDATA[3], posedge WCLK, 1.0);
   $setup(negedge WDATA[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[3], 1.0);
   $hold(posedge WCLK, negedge WDATA[3], 1.0);
   $setup(posedge WDATA[4], posedge WCLK, 1.0);
   $setup(negedge WDATA[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[4], 1.0);
   $hold(posedge WCLK, negedge WDATA[4], 1.0);
   $setup(posedge WDATA[5], posedge WCLK, 1.0);
   $setup(negedge WDATA[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[5], 1.0);
   $hold(posedge WCLK, negedge WDATA[5], 1.0);
   $setup(posedge WDATA[6], posedge WCLK, 1.0);
   $setup(negedge WDATA[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[6], 1.0);
   $hold(posedge WCLK, negedge WDATA[6], 1.0);
   $setup(posedge WDATA[7], posedge WCLK, 1.0);
   $setup(negedge WDATA[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[7], 1.0);
   $hold(posedge WCLK, negedge WDATA[7], 1.0);
   $setup(posedge WCLKE, posedge WCLK, 1.0);
   $setup(negedge WCLKE, posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WCLKE, 1.0);
   $hold(posedge WCLK, negedge WCLKE, 1.0);
   $setup(posedge WE, posedge WCLK, 1.0);
   $setup(negedge WE, posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WE, 1.0);
   $hold(posedge WCLK, negedge WE, 1.0);
   $setup(posedge RADDR[0], posedge RCLK, 1.0);
   $setup(negedge RADDR[0], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[0], 1.0);
   $hold(posedge RCLK, negedge RADDR[0], 1.0);
   $setup(posedge RADDR[1], posedge RCLK, 1.0);
   $setup(negedge RADDR[1], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[1], 1.0);
   $hold(posedge RCLK, negedge RADDR[1], 1.0);
   $setup(posedge RADDR[2], posedge RCLK, 1.0);
   $setup(negedge RADDR[2], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[2], 1.0);
   $hold(posedge RCLK, negedge RADDR[2], 1.0);
   $setup(posedge RADDR[3], posedge RCLK, 1.0);
   $setup(negedge RADDR[3], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[3], 1.0);
   $hold(posedge RCLK, negedge RADDR[3], 1.0);
   $setup(posedge RADDR[4], posedge RCLK, 1.0);
   $setup(negedge RADDR[4], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[4], 1.0);
   $hold(posedge RCLK, negedge RADDR[4], 1.0);
   $setup(posedge RADDR[5], posedge RCLK, 1.0);
   $setup(negedge RADDR[5], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[5], 1.0);
   $hold(posedge RCLK, negedge RADDR[5], 1.0);
   $setup(posedge RADDR[6], posedge RCLK, 1.0);
   $setup(negedge RADDR[6], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[6], 1.0);
   $hold(posedge RCLK, negedge RADDR[6], 1.0);
   $setup(posedge RADDR[7], posedge RCLK, 1.0);
   $setup(negedge RADDR[7], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[7], 1.0);
   $hold(posedge RCLK, negedge RADDR[7], 1.0);
   $setup(posedge RADDR[8], posedge RCLK, 1.0);
   $setup(negedge RADDR[8], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[8], 1.0);
   $hold(posedge RCLK, negedge RADDR[8], 1.0);
   $setup(posedge RCLKE, posedge RCLK, 1.0);
   $setup(negedge RCLKE, posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RCLKE, 1.0);
   $hold(posedge RCLK, negedge RCLKE, 1.0);
   $setup(posedge RE, posedge RCLK, 1.0);
   $setup(negedge RE, posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RE, 1.0);
   $hold(posedge RCLK, negedge RE, 1.0);

endspecify
`endif

endmodule //SB_RAM512x8


`timescale 1ps/1ps
module SB_RAM512x8NR (RDATA, RCLKN, RCLKE, RE, RADDR, WCLK, WCLKE, WE, WADDR, WDATA);
output [7:0] RDATA;
input RCLKN;
input RCLKE;
input RE;
input [8:0] RADDR;
input WCLK;
input WCLKE;
input WE;
input [8:0] WADDR;
input [7:0] WDATA;

parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

wire RCLK;
assign (weak0, weak1) RCLKE =1'b1 ;
assign (weak0, weak1) RE =1'b0 ;
assign (weak0, weak1) WCLKE =1'b1 ;
assign (weak0, weak1) WE =1'b0 ;
assign RCLK = ~RCLKN;

SB_RAM512x8 sb_ram512X8r_inst (
	.RDATA(RDATA),
	.RCLK(RCLK),
	.RCLKE(RCLKE),
	.RE(RE),
	.RADDR(RADDR),
	.WCLK(WCLK),
	.WCLKE(WCLKE),
	.WE(WE),
	.WADDR(WADDR),
	.WDATA(WDATA));

defparam sb_ram512X8r_inst.INIT_0 = INIT_0;
defparam sb_ram512X8r_inst.INIT_1 = INIT_1;
defparam sb_ram512X8r_inst.INIT_2 = INIT_2;
defparam sb_ram512X8r_inst.INIT_3 = INIT_3;
defparam sb_ram512X8r_inst.INIT_4 = INIT_4;
defparam sb_ram512X8r_inst.INIT_5 = INIT_5;
defparam sb_ram512X8r_inst.INIT_6 = INIT_6;
defparam sb_ram512X8r_inst.INIT_7 = INIT_7;
defparam sb_ram512X8r_inst.INIT_8 = INIT_8;
defparam sb_ram512X8r_inst.INIT_9 = INIT_9;
defparam sb_ram512X8r_inst.INIT_A = INIT_A;
defparam sb_ram512X8r_inst.INIT_B = INIT_B;
defparam sb_ram512X8r_inst.INIT_C = INIT_C;
defparam sb_ram512X8r_inst.INIT_D = INIT_D;
defparam sb_ram512X8r_inst.INIT_E = INIT_E;
defparam sb_ram512X8r_inst.INIT_F = INIT_F;

`ifdef TIMINGCHECK
specify
   (RCLKN *> RDATA[0]) = (1.0, 1.0);
   (RCLKN *> RDATA[1]) = (1.0, 1.0);
   (RCLKN *> RDATA[2]) = (1.0, 1.0);
   (RCLKN *> RDATA[3]) = (1.0, 1.0);
   (RCLKN *> RDATA[4]) = (1.0, 1.0);
   (RCLKN *> RDATA[5]) = (1.0, 1.0);
   (RCLKN *> RDATA[6]) = (1.0, 1.0);
   (RCLKN *> RDATA[7]) = (1.0, 1.0);
   $setup(posedge WADDR[0], posedge WCLK, 1.0);
   $setup(negedge WADDR[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[0], 1.0);
   $hold(posedge WCLK, negedge WADDR[0], 1.0);
   $setup(posedge WADDR[1], posedge WCLK, 1.0);
   $setup(negedge WADDR[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[1], 1.0);
   $hold(posedge WCLK, negedge WADDR[1], 1.0);
   $setup(posedge WADDR[2], posedge WCLK, 1.0);
   $setup(negedge WADDR[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[2], 1.0);
   $hold(posedge WCLK, negedge WADDR[2], 1.0);
   $setup(posedge WADDR[3], posedge WCLK, 1.0);
   $setup(negedge WADDR[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[3], 1.0);
   $hold(posedge WCLK, negedge WADDR[3], 1.0);
   $setup(posedge WADDR[4], posedge WCLK, 1.0);
   $setup(negedge WADDR[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[4], 1.0);
   $hold(posedge WCLK, negedge WADDR[4], 1.0);
   $setup(posedge WADDR[5], posedge WCLK, 1.0);
   $setup(negedge WADDR[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[5], 1.0);
   $hold(posedge WCLK, negedge WADDR[5], 1.0);
   $setup(posedge WADDR[6], posedge WCLK, 1.0);
   $setup(negedge WADDR[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[6], 1.0);
   $hold(posedge WCLK, negedge WADDR[6], 1.0);
   $setup(posedge WADDR[7], posedge WCLK, 1.0);
   $setup(negedge WADDR[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[7], 1.0);
   $hold(posedge WCLK, negedge WADDR[7], 1.0);
   $setup(posedge WADDR[8], posedge WCLK, 1.0);
   $setup(negedge WADDR[8], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[8], 1.0);
   $hold(posedge WCLK, negedge WADDR[8], 1.0);
   $setup(posedge WDATA[0], posedge WCLK, 1.0);
   $setup(negedge WDATA[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[0], 1.0);
   $hold(posedge WCLK, negedge WDATA[0], 1.0);
   $setup(posedge WDATA[1], posedge WCLK, 1.0);
   $setup(negedge WDATA[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[1], 1.0);
   $hold(posedge WCLK, negedge WDATA[1], 1.0);
   $setup(posedge WDATA[2], posedge WCLK, 1.0);
   $setup(negedge WDATA[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[2], 1.0);
   $hold(posedge WCLK, negedge WDATA[2], 1.0);
   $setup(posedge WDATA[3], posedge WCLK, 1.0);
   $setup(negedge WDATA[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[3], 1.0);
   $hold(posedge WCLK, negedge WDATA[3], 1.0);
   $setup(posedge WDATA[4], posedge WCLK, 1.0);
   $setup(negedge WDATA[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[4], 1.0);
   $hold(posedge WCLK, negedge WDATA[4], 1.0);
   $setup(posedge WDATA[5], posedge WCLK, 1.0);
   $setup(negedge WDATA[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[5], 1.0);
   $hold(posedge WCLK, negedge WDATA[5], 1.0);
   $setup(posedge WDATA[6], posedge WCLK, 1.0);
   $setup(negedge WDATA[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[6], 1.0);
   $hold(posedge WCLK, negedge WDATA[6], 1.0);
   $setup(posedge WDATA[7], posedge WCLK, 1.0);
   $setup(negedge WDATA[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[7], 1.0);
   $hold(posedge WCLK, negedge WDATA[7], 1.0);
   $setup(posedge WCLKE, posedge WCLK, 1.0);
   $setup(negedge WCLKE, posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WCLKE, 1.0);
   $hold(posedge WCLK, negedge WCLKE, 1.0);
   $setup(posedge WE, posedge WCLK, 1.0);
   $setup(negedge WE, posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WE, 1.0);
   $hold(posedge WCLK, negedge WE, 1.0);
   $setup(posedge RADDR[0], posedge RCLKN, 1.0);
   $setup(negedge RADDR[0], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[0], 1.0);
   $hold(posedge RCLKN, negedge RADDR[0], 1.0);
   $setup(posedge RADDR[1], posedge RCLKN, 1.0);
   $setup(negedge RADDR[1], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[1], 1.0);
   $hold(posedge RCLKN, negedge RADDR[1], 1.0);
   $setup(posedge RADDR[2], posedge RCLKN, 1.0);
   $setup(negedge RADDR[2], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[2], 1.0);
   $hold(posedge RCLKN, negedge RADDR[2], 1.0);
   $setup(posedge RADDR[3], posedge RCLKN, 1.0);
   $setup(negedge RADDR[3], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[3], 1.0);
   $hold(posedge RCLKN, negedge RADDR[3], 1.0);
   $setup(posedge RADDR[4], posedge RCLKN, 1.0);
   $setup(negedge RADDR[4], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[4], 1.0);
   $hold(posedge RCLKN, negedge RADDR[4], 1.0);
   $setup(posedge RADDR[5], posedge RCLKN, 1.0);
   $setup(negedge RADDR[5], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[5], 1.0);
   $hold(posedge RCLKN, negedge RADDR[5], 1.0);
   $setup(posedge RADDR[6], posedge RCLKN, 1.0);
   $setup(negedge RADDR[6], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[6], 1.0);
   $hold(posedge RCLKN, negedge RADDR[6], 1.0);
   $setup(posedge RADDR[7], posedge RCLKN, 1.0);
   $setup(negedge RADDR[7], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[7], 1.0);
   $hold(posedge RCLKN, negedge RADDR[7], 1.0);
   $setup(posedge RADDR[8], posedge RCLKN, 1.0);
   $setup(negedge RADDR[8], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[8], 1.0);
   $hold(posedge RCLKN, negedge RADDR[8], 1.0);
   $setup(posedge RCLKE, posedge RCLKN, 1.0);
   $setup(negedge RCLKE, posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RCLKE, 1.0);
   $hold(posedge RCLKN, negedge RCLKE, 1.0);
   $setup(posedge RE, posedge RCLKN, 1.0);
   $setup(negedge RE, posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RE, 1.0);
   $hold(posedge RCLKN, negedge RE, 1.0);
   $recovery(posedge RCLKN, posedge WCLK, 1.0);
   $recovery(negedge RCLKN, posedge WCLK, 1.0);
   $removal(posedge RCLKN, posedge WCLK, 1.0);
   $removal(negedge RCLKN, posedge WCLK, 1.0);
   $recovery(posedge WCLK, posedge RCLKN, 1.0);
   $recovery(negedge WCLK, posedge RCLKN, 1.0);
   $removal(posedge WCLK, posedge RCLKN, 1.0);
   $removal(negedge WCLK, posedge RCLKN, 1.0);

endspecify
`endif
endmodule //SB_RAM512x8NR


`timescale 1ps/1ps
module SB_RAM512x8NW (RDATA, RCLK, RCLKE, RE, RADDR, WCLKN, WCLKE, WE, WADDR, WDATA);
output [7:0] RDATA;
input RCLK;
input RCLKE;
input RE;
input [8:0] RADDR;
input WCLKN;
input WCLKE;
input WE;
input [8:0] WADDR;
input [7:0] WDATA;

parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

wire WCLK;
assign (weak0, weak1) RCLKE =1'b1 ;
assign (weak0, weak1) RE =1'b0 ;
assign (weak0, weak1) WCLKE =1'b1 ;
assign (weak0, weak1) WE =1'b0 ;
assign WCLK = ~WCLKN;

SB_RAM512x8 sb_ram512X8w_inst (
	.RDATA(RDATA),
	.RCLK(RCLK),
	.RCLKE(RCLKE),
	.RE(RE),
	.RADDR(RADDR),
	.WCLK(WCLK),
	.WCLKE(WCLKE),
	.WE(WE),
	.WADDR(WADDR),
	.WDATA(WDATA));

defparam sb_ram512X8w_inst.INIT_0 = INIT_0;
defparam sb_ram512X8w_inst.INIT_1 = INIT_1;
defparam sb_ram512X8w_inst.INIT_2 = INIT_2;
defparam sb_ram512X8w_inst.INIT_3 = INIT_3;
defparam sb_ram512X8w_inst.INIT_4 = INIT_4;
defparam sb_ram512X8w_inst.INIT_5 = INIT_5;
defparam sb_ram512X8w_inst.INIT_6 = INIT_6;
defparam sb_ram512X8w_inst.INIT_7 = INIT_7;
defparam sb_ram512X8w_inst.INIT_8 = INIT_8;
defparam sb_ram512X8w_inst.INIT_9 = INIT_9;
defparam sb_ram512X8w_inst.INIT_A = INIT_A;
defparam sb_ram512X8w_inst.INIT_B = INIT_B;
defparam sb_ram512X8w_inst.INIT_C = INIT_C;
defparam sb_ram512X8w_inst.INIT_D = INIT_D;
defparam sb_ram512X8w_inst.INIT_E = INIT_E;
defparam sb_ram512X8w_inst.INIT_F = INIT_F;

`ifdef TIMINGCHECK
specify
   (RCLK *> RDATA[0]) = (1.0, 1.0);
   (RCLK *> RDATA[1]) = (1.0, 1.0);
   (RCLK *> RDATA[2]) = (1.0, 1.0);
   (RCLK *> RDATA[3]) = (1.0, 1.0);
   (RCLK *> RDATA[4]) = (1.0, 1.0);
   (RCLK *> RDATA[5]) = (1.0, 1.0);
   (RCLK *> RDATA[6]) = (1.0, 1.0);
   (RCLK *> RDATA[7]) = (1.0, 1.0);
   $setup(posedge WADDR[0], posedge WCLKN, 1.0);
   $setup(negedge WADDR[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[0], 1.0);
   $hold(posedge WCLKN, negedge WADDR[0], 1.0);
   $setup(posedge WADDR[1], posedge WCLKN, 1.0);
   $setup(negedge WADDR[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[1], 1.0);
   $hold(posedge WCLKN, negedge WADDR[1], 1.0);
   $setup(posedge WADDR[2], posedge WCLKN, 1.0);
   $setup(negedge WADDR[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[2], 1.0);
   $hold(posedge WCLKN, negedge WADDR[2], 1.0);
   $setup(posedge WADDR[3], posedge WCLKN, 1.0);
   $setup(negedge WADDR[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[3], 1.0);
   $hold(posedge WCLKN, negedge WADDR[3], 1.0);
   $setup(posedge WADDR[4], posedge WCLKN, 1.0);
   $setup(negedge WADDR[4], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[4], 1.0);
   $hold(posedge WCLKN, negedge WADDR[4], 1.0);
   $setup(posedge WADDR[5], posedge WCLKN, 1.0);
   $setup(negedge WADDR[5], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[5], 1.0);
   $hold(posedge WCLKN, negedge WADDR[5], 1.0);
   $setup(posedge WADDR[6], posedge WCLKN, 1.0);
   $setup(negedge WADDR[6], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[6], 1.0);
   $hold(posedge WCLKN, negedge WADDR[6], 1.0);
   $setup(posedge WADDR[7], posedge WCLKN, 1.0);
   $setup(negedge WADDR[7], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[7], 1.0);
   $hold(posedge WCLKN, negedge WADDR[7], 1.0);
   $setup(posedge WADDR[8], posedge WCLKN, 1.0);
   $setup(negedge WADDR[8], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[8], 1.0);
   $hold(posedge WCLKN, negedge WADDR[8], 1.0);
   $setup(posedge WDATA[0], posedge WCLKN, 1.0);
   $setup(negedge WDATA[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[0], 1.0);
   $hold(posedge WCLKN, negedge WDATA[0], 1.0);
   $setup(posedge WDATA[1], posedge WCLKN, 1.0);
   $setup(negedge WDATA[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[1], 1.0);
   $hold(posedge WCLKN, negedge WDATA[1], 1.0);
   $setup(posedge WDATA[2], posedge WCLKN, 1.0);
   $setup(negedge WDATA[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[2], 1.0);
   $hold(posedge WCLKN, negedge WDATA[2], 1.0);
   $setup(posedge WDATA[3], posedge WCLKN, 1.0);
   $setup(negedge WDATA[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[3], 1.0);
   $hold(posedge WCLKN, negedge WDATA[3], 1.0);
   $setup(posedge WDATA[4], posedge WCLKN, 1.0);
   $setup(negedge WDATA[4], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[4], 1.0);
   $hold(posedge WCLKN, negedge WDATA[4], 1.0);
   $setup(posedge WDATA[5], posedge WCLKN, 1.0);
   $setup(negedge WDATA[5], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[5], 1.0);
   $hold(posedge WCLKN, negedge WDATA[5], 1.0);
   $setup(posedge WDATA[6], posedge WCLKN, 1.0);
   $setup(negedge WDATA[6], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[6], 1.0);
   $hold(posedge WCLKN, negedge WDATA[6], 1.0);
   $setup(posedge WDATA[7], posedge WCLKN, 1.0);
   $setup(negedge WDATA[7], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[7], 1.0);
   $hold(posedge WCLKN, negedge WDATA[7], 1.0);
   $setup(posedge WCLKE, posedge WCLKN, 1.0);
   $setup(negedge WCLKE, posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WCLKE, 1.0);
   $hold(posedge WCLKN, negedge WCLKE, 1.0);
   $setup(posedge WE, posedge WCLKN, 1.0);
   $setup(negedge WE, posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WE, 1.0);
   $hold(posedge WCLKN, negedge WE, 1.0);
   $setup(posedge RADDR[0], posedge RCLK, 1.0);
   $setup(negedge RADDR[0], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[0], 1.0);
   $hold(posedge RCLK, negedge RADDR[0], 1.0);
   $setup(posedge RADDR[1], posedge RCLK, 1.0);
   $setup(negedge RADDR[1], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[1], 1.0);
   $hold(posedge RCLK, negedge RADDR[1], 1.0);
   $setup(posedge RADDR[2], posedge RCLK, 1.0);
   $setup(negedge RADDR[2], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[2], 1.0);
   $hold(posedge RCLK, negedge RADDR[2], 1.0);
   $setup(posedge RADDR[3], posedge RCLK, 1.0);
   $setup(negedge RADDR[3], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[3], 1.0);
   $hold(posedge RCLK, negedge RADDR[3], 1.0);
   $setup(posedge RADDR[4], posedge RCLK, 1.0);
   $setup(negedge RADDR[4], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[4], 1.0);
   $hold(posedge RCLK, negedge RADDR[4], 1.0);
   $setup(posedge RADDR[5], posedge RCLK, 1.0);
   $setup(negedge RADDR[5], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[5], 1.0);
   $hold(posedge RCLK, negedge RADDR[5], 1.0);
   $setup(posedge RADDR[6], posedge RCLK, 1.0);
   $setup(negedge RADDR[6], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[6], 1.0);
   $hold(posedge RCLK, negedge RADDR[6], 1.0);
   $setup(posedge RADDR[7], posedge RCLK, 1.0);
   $setup(negedge RADDR[7], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[7], 1.0);
   $hold(posedge RCLK, negedge RADDR[7], 1.0);
   $setup(posedge RADDR[8], posedge RCLK, 1.0);
   $setup(negedge RADDR[8], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[8], 1.0);
   $hold(posedge RCLK, negedge RADDR[8], 1.0);
   $setup(posedge RCLKE, posedge RCLK, 1.0);
   $setup(negedge RCLKE, posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RCLKE, 1.0);
   $hold(posedge RCLK, negedge RCLKE, 1.0);
   $setup(posedge RE, posedge RCLK, 1.0);
   $setup(negedge RE, posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RE, 1.0);
   $hold(posedge RCLK, negedge RE, 1.0);
   $recovery(posedge RCLK, posedge WCLKN, 1.0);
   $recovery(negedge RCLK, posedge WCLKN, 1.0);
   $removal(posedge RCLK, posedge WCLKN, 1.0);
   $removal(negedge RCLK, posedge WCLKN, 1.0);
   $recovery(posedge WCLKN, posedge RCLK, 1.0);
   $recovery(negedge WCLKN, posedge RCLK, 1.0);
   $removal(posedge WCLKN, posedge RCLK, 1.0);
   $removal(negedge WCLKN, posedge RCLK, 1.0);

endspecify
`endif
endmodule //SB_RAM512x8NW


`timescale 1ps/1ps
module SB_RAM512x8NRNW (RDATA, RCLKN, RCLKE, RE, RADDR, WCLKN, WCLKE, WE, WADDR, WDATA);
output [7:0] RDATA;
input RCLKN;
input RCLKE;
input RE;
input [8:0] RADDR;
input WCLKN;
input WCLKE;
input WE;
input [8:0] WADDR;
input [7:0] WDATA;

parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

wire RCLK, WCLK;
assign (weak0, weak1) RCLKE =1'b1 ;
assign (weak0, weak1) RE =1'b0 ;
assign (weak0, weak1) WCLKE =1'b1 ;
assign (weak0, weak1) WE =1'b0 ;
assign RCLK = ~RCLKN;
assign WCLK = ~WCLKN;

SB_RAM512x8 sb_ram512X8rw_inst (
	.RDATA(RDATA),
	.RCLK(RCLK),
	.RCLKE(RCLKE),
	.RE(RE),
	.RADDR(RADDR),
	.WCLK(WCLK),
	.WCLKE(WCLKE),
	.WE(WE),
	.WADDR(WADDR),
	.WDATA(WDATA));

defparam sb_ram512X8rw_inst.INIT_0 = INIT_0;
defparam sb_ram512X8rw_inst.INIT_1 = INIT_1;
defparam sb_ram512X8rw_inst.INIT_2 = INIT_2;
defparam sb_ram512X8rw_inst.INIT_3 = INIT_3;
defparam sb_ram512X8rw_inst.INIT_4 = INIT_4;
defparam sb_ram512X8rw_inst.INIT_5 = INIT_5;
defparam sb_ram512X8rw_inst.INIT_6 = INIT_6;
defparam sb_ram512X8rw_inst.INIT_7 = INIT_7;
defparam sb_ram512X8rw_inst.INIT_8 = INIT_8;
defparam sb_ram512X8rw_inst.INIT_9 = INIT_9;
defparam sb_ram512X8rw_inst.INIT_A = INIT_A;
defparam sb_ram512X8rw_inst.INIT_B = INIT_B;
defparam sb_ram512X8rw_inst.INIT_C = INIT_C;
defparam sb_ram512X8rw_inst.INIT_D = INIT_D;
defparam sb_ram512X8rw_inst.INIT_E = INIT_E;
defparam sb_ram512X8rw_inst.INIT_F = INIT_F;

`ifdef TIMINGCHECK
specify
   (RCLKN *> RDATA[0]) = (1.0, 1.0);
   (RCLKN *> RDATA[1]) = (1.0, 1.0);
   (RCLKN *> RDATA[2]) = (1.0, 1.0);
   (RCLKN *> RDATA[3]) = (1.0, 1.0);
   (RCLKN *> RDATA[4]) = (1.0, 1.0);
   (RCLKN *> RDATA[5]) = (1.0, 1.0);
   (RCLKN *> RDATA[6]) = (1.0, 1.0);
   (RCLKN *> RDATA[7]) = (1.0, 1.0);
   $setup(posedge WADDR[0], posedge WCLKN, 1.0);
   $setup(negedge WADDR[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[0], 1.0);
   $hold(posedge WCLKN, negedge WADDR[0], 1.0);
   $setup(posedge WADDR[1], posedge WCLKN, 1.0);
   $setup(negedge WADDR[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[1], 1.0);
   $hold(posedge WCLKN, negedge WADDR[1], 1.0);
   $setup(posedge WADDR[2], posedge WCLKN, 1.0);
   $setup(negedge WADDR[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[2], 1.0);
   $hold(posedge WCLKN, negedge WADDR[2], 1.0);
   $setup(posedge WADDR[3], posedge WCLKN, 1.0);
   $setup(negedge WADDR[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[3], 1.0);
   $hold(posedge WCLKN, negedge WADDR[3], 1.0);
   $setup(posedge WADDR[4], posedge WCLKN, 1.0);
   $setup(negedge WADDR[4], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[4], 1.0);
   $hold(posedge WCLKN, negedge WADDR[4], 1.0);
   $setup(posedge WADDR[5], posedge WCLKN, 1.0);
   $setup(negedge WADDR[5], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[5], 1.0);
   $hold(posedge WCLKN, negedge WADDR[5], 1.0);
   $setup(posedge WADDR[6], posedge WCLKN, 1.0);
   $setup(negedge WADDR[6], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[6], 1.0);
   $hold(posedge WCLKN, negedge WADDR[6], 1.0);
   $setup(posedge WADDR[7], posedge WCLKN, 1.0);
   $setup(negedge WADDR[7], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[7], 1.0);
   $hold(posedge WCLKN, negedge WADDR[7], 1.0);
   $setup(posedge WADDR[8], posedge WCLKN, 1.0);
   $setup(negedge WADDR[8], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[8], 1.0);
   $hold(posedge WCLKN, negedge WADDR[8], 1.0);
   $setup(posedge WDATA[0], posedge WCLKN, 1.0);
   $setup(negedge WDATA[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[0], 1.0);
   $hold(posedge WCLKN, negedge WDATA[0], 1.0);
   $setup(posedge WDATA[1], posedge WCLKN, 1.0);
   $setup(negedge WDATA[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[1], 1.0);
   $hold(posedge WCLKN, negedge WDATA[1], 1.0);
   $setup(posedge WDATA[2], posedge WCLKN, 1.0);
   $setup(negedge WDATA[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[2], 1.0);
   $hold(posedge WCLKN, negedge WDATA[2], 1.0);
   $setup(posedge WDATA[3], posedge WCLKN, 1.0);
   $setup(negedge WDATA[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[3], 1.0);
   $hold(posedge WCLKN, negedge WDATA[3], 1.0);
   $setup(posedge WDATA[4], posedge WCLKN, 1.0);
   $setup(negedge WDATA[4], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[4], 1.0);
   $hold(posedge WCLKN, negedge WDATA[4], 1.0);
   $setup(posedge WDATA[5], posedge WCLKN, 1.0);
   $setup(negedge WDATA[5], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[5], 1.0);
   $hold(posedge WCLKN, negedge WDATA[5], 1.0);
   $setup(posedge WDATA[6], posedge WCLKN, 1.0);
   $setup(negedge WDATA[6], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[6], 1.0);
   $hold(posedge WCLKN, negedge WDATA[6], 1.0);
   $setup(posedge WDATA[7], posedge WCLKN, 1.0);
   $setup(negedge WDATA[7], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[7], 1.0);
   $hold(posedge WCLKN, negedge WDATA[7], 1.0);
   $setup(posedge WCLKE, posedge WCLKN, 1.0);
   $setup(negedge WCLKE, posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WCLKE, 1.0);
   $hold(posedge WCLKN, negedge WCLKE, 1.0);
   $setup(posedge WE, posedge WCLKN, 1.0);
   $setup(negedge WE, posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WE, 1.0);
   $hold(posedge WCLKN, negedge WE, 1.0);
   $setup(posedge RADDR[0], posedge RCLKN, 1.0);
   $setup(negedge RADDR[0], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[0], 1.0);
   $hold(posedge RCLKN, negedge RADDR[0], 1.0);
   $setup(posedge RADDR[1], posedge RCLKN, 1.0);
   $setup(negedge RADDR[1], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[1], 1.0);
   $hold(posedge RCLKN, negedge RADDR[1], 1.0);
   $setup(posedge RADDR[2], posedge RCLKN, 1.0);
   $setup(negedge RADDR[2], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[2], 1.0);
   $hold(posedge RCLKN, negedge RADDR[2], 1.0);
   $setup(posedge RADDR[3], posedge RCLKN, 1.0);
   $setup(negedge RADDR[3], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[3], 1.0);
   $hold(posedge RCLKN, negedge RADDR[3], 1.0);
   $setup(posedge RADDR[4], posedge RCLKN, 1.0);
   $setup(negedge RADDR[4], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[4], 1.0);
   $hold(posedge RCLKN, negedge RADDR[4], 1.0);
   $setup(posedge RADDR[5], posedge RCLKN, 1.0);
   $setup(negedge RADDR[5], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[5], 1.0);
   $hold(posedge RCLKN, negedge RADDR[5], 1.0);
   $setup(posedge RADDR[6], posedge RCLKN, 1.0);
   $setup(negedge RADDR[6], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[6], 1.0);
   $hold(posedge RCLKN, negedge RADDR[6], 1.0);
   $setup(posedge RADDR[7], posedge RCLKN, 1.0);
   $setup(negedge RADDR[7], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[7], 1.0);
   $hold(posedge RCLKN, negedge RADDR[7], 1.0);
   $setup(posedge RADDR[8], posedge RCLKN, 1.0);
   $setup(negedge RADDR[8], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[8], 1.0);
   $hold(posedge RCLKN, negedge RADDR[8], 1.0);
   $setup(posedge RCLKE, posedge RCLKN, 1.0);
   $setup(negedge RCLKE, posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RCLKE, 1.0);
   $hold(posedge RCLKN, negedge RCLKE, 1.0);
   $setup(posedge RE, posedge RCLKN, 1.0);
   $setup(negedge RE, posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RE, 1.0);
   $hold(posedge RCLKN, negedge RE, 1.0);
   $recovery(posedge RCLKN, posedge WCLKN, 1.0);
   $recovery(negedge RCLKN, posedge WCLKN, 1.0);
   $removal(posedge RCLKN, posedge WCLKN, 1.0);
   $removal(negedge RCLKN, posedge WCLKN, 1.0);
   $recovery(posedge WCLKN, posedge RCLKN, 1.0);
   $recovery(negedge WCLKN, posedge RCLKN, 1.0);
   $removal(posedge WCLKN, posedge RCLKN, 1.0);
   $removal(negedge WCLKN, posedge RCLKN, 1.0);

endspecify
`endif
endmodule //SB_RAM512x8NRNW


`timescale 1ps/1ps
module SB_RAM1024x4 (RDATA, RCLK, RCLKE, RE, RADDR, WCLK, WCLKE, WE, WADDR, WDATA);
output [3:0] RDATA;
input RCLK;
input RCLKE;
input RE;
input [9:0] RADDR;
input WCLK;
input WCLKE;
input WE;
input [9:0] WADDR;
input [3:0] WDATA;

parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

// local Parameters
localparam			CLOCK_PERIOD = 200;	//
localparam 			DELAY	= (CLOCK_PERIOD/10);		// Clock-to-output delay. Zero
							// time delays can be confusing
							// and sometimes cause problems.
localparam 			BUS_WIDTH = 4;		// Width of RAM (number of bits)

localparam 			ADDRESS_BUS_SIZE = 10;	// Number of bits required to
							// represent the RAM address

localparam   ADDRESSABLE_SPACE  = 2**ADDRESS_BUS_SIZE;	// Decimal address range [2^Size:0]


// SIGNAL DECLARATIONS
wire			   	WCLK_g, RCLK_g;
reg 				WCLKE_sync, RCLKE_sync; 
assign (weak0, weak1) RCLKE =1'b1 ;
assign (weak0, weak1) RE =1'b0 ;
assign (weak0, weak1) WCLKE =1'b1 ;
assign (weak0, weak1) WE =1'b0 ;
reg	Memory	[BUS_WIDTH*ADDRESSABLE_SPACE-1:0];
// 
event Read_e, Write_e;

//////////////////// Collision detect begins here ///////////////////////////////
localparam 	TRUE = 1'b1;
localparam	FALSE = 1'b0;
reg 		Time_Collision_Detected = 1'b0;
wire		Address_Collision_Detected;

event Collision_e;

time COLLISION_TIME_WINDOW = (CLOCK_PERIOD/8); // This is an arbitray value, but is better than using an absolute 
						    // value, because the actual time window depends on the actual silicon 
						    // implementation. Thus the test is indicative of an Error and not
						    // guaranteed to be an error. Even so this is usefull.
time time_WCLK_RCLK, time_WCLK, time_RCLK;


//function reg Check_Timed_Window_Violation;
function	Check_Timed_Window_Violation;	//	by Jeffrey
input T1, T2, Minimum_Time_Window;
time T1, T2;
time Minimum_Time_Window;
time Difference;	
	begin
		Difference = (T1 - T2);
		if (Difference < 0) Difference = -Difference;
		Check_Timed_Window_Violation = (Difference < Minimum_Time_Window);
	end
endfunction


initial begin
       time_WCLK = CLOCK_PERIOD;	// Arbitrary initialisation value, ensure no window collison error on first clock edge.
       time_RCLK = (CLOCK_PERIOD*8);	// Arbitrary initialisation difference value, ensure no collision error on first clock edge.					
end

integer	i,j;


initial	//	initialize ram_4k by parameter, section by section
begin
	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[BUS_WIDTH*i+j]	=	INIT_0[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*1+BUS_WIDTH*i+j]	=	INIT_1[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*2+BUS_WIDTH*i+j]	=	INIT_2[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*3+BUS_WIDTH*i+j]	=	INIT_3[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*4+BUS_WIDTH*i+j]	=	INIT_4[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*5+BUS_WIDTH*i+j]	=	INIT_5[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*6+BUS_WIDTH*i+j]	=	INIT_6[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*7+BUS_WIDTH*i+j]	=	INIT_7[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*8+BUS_WIDTH*i+j]	=	INIT_8[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*9+BUS_WIDTH*i+j]	=	INIT_9[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*10+BUS_WIDTH*i+j]	=	INIT_A[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*11+BUS_WIDTH*i+j]	=	INIT_B[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*12+BUS_WIDTH*i+j]	=	INIT_C[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*13+BUS_WIDTH*i+j]	=	INIT_D[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*14+BUS_WIDTH*i+j]	=	INIT_E[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*15+BUS_WIDTH*i+j]	=	INIT_F[BUS_WIDTH*i+j];
	end

end

assign Address_Collision_Detected = ((RE & WE & WCLKE & RCLKE)&(WADDR == RADDR)); 


always @(WCLK or WCLKE) 
begin 
	if(~WCLK)
	WCLKE_sync = WCLKE;   	
end 

always @(RCLK or RCLKE) 
begin 
	if (~RCLK)
	RCLKE_sync = RCLKE; 	
end 

assign WCLK_g = WCLK & WCLKE_sync;
assign RCLK_g = RCLK & RCLKE_sync;

always @(posedge WCLK_g) begin
	time_WCLK = $time;
end

always @(posedge RCLK_g) begin
    	time_RCLK = $time;
end
integer	SB_RAM1024X4_RDATA_log_file;					//.....................
initial	SB_RAM1024X4_RDATA_log_file=("SB_RAM1024X4_RDATA_log_file.txt");	//.....................
always @(posedge WCLK_g) begin

	Time_Collision_Detected = Check_Timed_Window_Violation(time_WCLK,time_RCLK,COLLISION_TIME_WINDOW);
        if (Time_Collision_Detected & Address_Collision_Detected)begin
        	$display("Warning: Write-Read collision detected, Data read value is X\n");
 		$display("WCLK Time: %.3f   RCLK Time:%.3f  ",time_WCLK, time_RCLK,"WADDR: %d   RADDR:%d\n",WADDR, RADDR); 
 		$fdisplay(SB_RAM1024X4_RDATA_log_file,"Warning: Write-Read collision detected, Data read value is X\n");
		$fdisplay(SB_RAM1024X4_RDATA_log_file,"WCLK Time: %.3f   RCLK Time:%.3f  ",time_WCLK, time_RCLK, "WADDR: %d   RADDR:%d\n",WADDR, RADDR); 	
 		-> Collision_e;
	end
end




//	code modify for universal verilog compiler

always @ (posedge WCLK_g)
begin
	if	(WE)
	begin
		-> Write_e;
		for	(i=0;i<=BUS_WIDTH-1; i=i+1)
		begin
			Memory[WADDR*BUS_WIDTH+i]	<=	WDATA[i];
		end
	end
end

//reg	[3:0]	RDATA = 0;
reg	[3:0]	RDATA;

initial
begin
   RDATA = $random;
end

// Look at the rising edge of the clock

always @ (posedge RCLK_g)
begin
	if	(RE)
	begin
		-> Read_e;
		if	(Time_Collision_Detected & Address_Collision_Detected) 
			RDATA <= 4'hX;
		else
			for	(i=0;i<=BUS_WIDTH-1;i=i+1)
				RDATA[i]	<= Memory[RADDR*BUS_WIDTH+i];
	end
end

`ifdef TIMINGCHECK
specify
   (RCLK *> RDATA[0]) = (1.0, 1.0);
   (RCLK *> RDATA[1]) = (1.0, 1.0);
   (RCLK *> RDATA[2]) = (1.0, 1.0);
   (RCLK *> RDATA[3]) = (1.0, 1.0);
   $setup(posedge WADDR[0], posedge WCLK, 1.0);
   $setup(negedge WADDR[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[0], 1.0);
   $hold(posedge WCLK, negedge WADDR[0], 1.0);
   $setup(posedge WADDR[1], posedge WCLK, 1.0);
   $setup(negedge WADDR[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[1], 1.0);
   $hold(posedge WCLK, negedge WADDR[1], 1.0);
   $setup(posedge WADDR[2], posedge WCLK, 1.0);
   $setup(negedge WADDR[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[2], 1.0);
   $hold(posedge WCLK, negedge WADDR[2], 1.0);
   $setup(posedge WADDR[3], posedge WCLK, 1.0);
   $setup(negedge WADDR[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[3], 1.0);
   $hold(posedge WCLK, negedge WADDR[3], 1.0);
   $setup(posedge WADDR[4], posedge WCLK, 1.0);
   $setup(negedge WADDR[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[4], 1.0);
   $hold(posedge WCLK, negedge WADDR[4], 1.0);
   $setup(posedge WADDR[5], posedge WCLK, 1.0);
   $setup(negedge WADDR[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[5], 1.0);
   $hold(posedge WCLK, negedge WADDR[5], 1.0);
   $setup(posedge WADDR[6], posedge WCLK, 1.0);
   $setup(negedge WADDR[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[6], 1.0);
   $hold(posedge WCLK, negedge WADDR[6], 1.0);
   $setup(posedge WADDR[7], posedge WCLK, 1.0);
   $setup(negedge WADDR[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[7], 1.0);
   $hold(posedge WCLK, negedge WADDR[7], 1.0);
   $setup(posedge WADDR[8], posedge WCLK, 1.0);
   $setup(negedge WADDR[8], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[8], 1.0);
   $hold(posedge WCLK, negedge WADDR[8], 1.0);
   $setup(posedge WADDR[9], posedge WCLK, 1.0);
   $setup(negedge WADDR[9], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[9], 1.0);
   $hold(posedge WCLK, negedge WADDR[9], 1.0);
   $setup(posedge WDATA[0], posedge WCLK, 1.0);
   $setup(negedge WDATA[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[0], 1.0);
   $hold(posedge WCLK, negedge WDATA[0], 1.0);
   $setup(posedge WDATA[1], posedge WCLK, 1.0);
   $setup(negedge WDATA[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[1], 1.0);
   $hold(posedge WCLK, negedge WDATA[1], 1.0);
   $setup(posedge WDATA[2], posedge WCLK, 1.0);
   $setup(negedge WDATA[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[2], 1.0);
   $hold(posedge WCLK, negedge WDATA[2], 1.0);
   $setup(posedge WDATA[3], posedge WCLK, 1.0);
   $setup(negedge WDATA[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[3], 1.0);
   $hold(posedge WCLK, negedge WDATA[3], 1.0);
   $setup(posedge WCLKE, posedge WCLK, 1.0);
   $setup(negedge WCLKE, posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WCLKE, 1.0);
   $hold(posedge WCLK, negedge WCLKE, 1.0);
   $setup(posedge WE, posedge WCLK, 1.0);
   $setup(negedge WE, posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WE, 1.0);
   $hold(posedge WCLK, negedge WE, 1.0);
   $setup(posedge RADDR[0], posedge RCLK, 1.0);
   $setup(negedge RADDR[0], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[0], 1.0);
   $hold(posedge RCLK, negedge RADDR[0], 1.0);
   $setup(posedge RADDR[1], posedge RCLK, 1.0);
   $setup(negedge RADDR[1], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[1], 1.0);
   $hold(posedge RCLK, negedge RADDR[1], 1.0);
   $setup(posedge RADDR[2], posedge RCLK, 1.0);
   $setup(negedge RADDR[2], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[2], 1.0);
   $hold(posedge RCLK, negedge RADDR[2], 1.0);
   $setup(posedge RADDR[3], posedge RCLK, 1.0);
   $setup(negedge RADDR[3], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[3], 1.0);
   $hold(posedge RCLK, negedge RADDR[3], 1.0);
   $setup(posedge RADDR[4], posedge RCLK, 1.0);
   $setup(negedge RADDR[4], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[4], 1.0);
   $hold(posedge RCLK, negedge RADDR[4], 1.0);
   $setup(posedge RADDR[5], posedge RCLK, 1.0);
   $setup(negedge RADDR[5], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[5], 1.0);
   $hold(posedge RCLK, negedge RADDR[5], 1.0);
   $setup(posedge RADDR[6], posedge RCLK, 1.0);
   $setup(negedge RADDR[6], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[6], 1.0);
   $hold(posedge RCLK, negedge RADDR[6], 1.0);
   $setup(posedge RADDR[7], posedge RCLK, 1.0);
   $setup(negedge RADDR[7], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[7], 1.0);
   $hold(posedge RCLK, negedge RADDR[7], 1.0);
   $setup(posedge RADDR[8], posedge RCLK, 1.0);
   $setup(negedge RADDR[8], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[8], 1.0);
   $hold(posedge RCLK, negedge RADDR[8], 1.0);
   $setup(posedge RADDR[9], posedge RCLK, 1.0);
   $setup(negedge RADDR[9], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[9], 1.0);
   $hold(posedge RCLK, negedge RADDR[9], 1.0);
   $setup(posedge RCLKE, posedge RCLK, 1.0);
   $setup(negedge RCLKE, posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RCLKE, 1.0);
   $hold(posedge RCLK, negedge RCLKE, 1.0);
   $setup(posedge RE, posedge RCLK, 1.0);
   $setup(negedge RE, posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RE, 1.0);
   $hold(posedge RCLK, negedge RE, 1.0);

endspecify
`endif


endmodule //SB_RAM1024x4


`timescale 1ps/1ps
module SB_RAM1024x4NR (RDATA, RCLKN, RCLKE, RE, RADDR, WCLK, WCLKE, WE, WADDR, WDATA);
output [3:0] RDATA;
input RCLKN;
input RCLKE;
input RE;
input [9:0] RADDR;
input WCLK;
input WCLKE;
input WE;
input [9:0] WADDR;
input [3:0] WDATA;

parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;


wire RCLK;
assign (weak0, weak1) RCLKE =1'b1 ;
assign (weak0, weak1) RE =1'b0 ;
assign (weak0, weak1) WCLKE =1'b1 ;
assign (weak0, weak1) WE =1'b0 ;
assign RCLK = ~RCLKN;

SB_RAM1024x4 sb_ram1024X4r_inst (
	.RDATA(RDATA),
	.RCLK(RCLK),
	.RCLKE(RCLKE),
	.RE(RE),
	.RADDR(RADDR),
	.WCLK(WCLK),
	.WCLKE(WCLKE),
	.WE(WE),
	.WADDR(WADDR),
	.WDATA(WDATA));

defparam sb_ram1024X4r_inst.INIT_0 = INIT_0;
defparam sb_ram1024X4r_inst.INIT_1 = INIT_1;
defparam sb_ram1024X4r_inst.INIT_2 = INIT_2;
defparam sb_ram1024X4r_inst.INIT_3 = INIT_3;
defparam sb_ram1024X4r_inst.INIT_4 = INIT_4;
defparam sb_ram1024X4r_inst.INIT_5 = INIT_5;
defparam sb_ram1024X4r_inst.INIT_6 = INIT_6;
defparam sb_ram1024X4r_inst.INIT_7 = INIT_7;
defparam sb_ram1024X4r_inst.INIT_8 = INIT_8;
defparam sb_ram1024X4r_inst.INIT_9 = INIT_9;
defparam sb_ram1024X4r_inst.INIT_A = INIT_A;
defparam sb_ram1024X4r_inst.INIT_B = INIT_B;
defparam sb_ram1024X4r_inst.INIT_C = INIT_C;
defparam sb_ram1024X4r_inst.INIT_D = INIT_D;
defparam sb_ram1024X4r_inst.INIT_E = INIT_E;
defparam sb_ram1024X4r_inst.INIT_F = INIT_F;

`ifdef TIMINGCHECK
specify
   (RCLKN *> RDATA[0]) = (1.0, 1.0);
   (RCLKN *> RDATA[1]) = (1.0, 1.0);
   (RCLKN *> RDATA[2]) = (1.0, 1.0);
   (RCLKN *> RDATA[3]) = (1.0, 1.0);
   $setup(posedge WADDR[0], posedge WCLK, 1.0);
   $setup(negedge WADDR[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[0], 1.0);
   $hold(posedge WCLK, negedge WADDR[0], 1.0);
   $setup(posedge WADDR[1], posedge WCLK, 1.0);
   $setup(negedge WADDR[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[1], 1.0);
   $hold(posedge WCLK, negedge WADDR[1], 1.0);
   $setup(posedge WADDR[2], posedge WCLK, 1.0);
   $setup(negedge WADDR[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[2], 1.0);
   $hold(posedge WCLK, negedge WADDR[2], 1.0);
   $setup(posedge WADDR[3], posedge WCLK, 1.0);
   $setup(negedge WADDR[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[3], 1.0);
   $hold(posedge WCLK, negedge WADDR[3], 1.0);
   $setup(posedge WADDR[4], posedge WCLK, 1.0);
   $setup(negedge WADDR[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[4], 1.0);
   $hold(posedge WCLK, negedge WADDR[4], 1.0);
   $setup(posedge WADDR[5], posedge WCLK, 1.0);
   $setup(negedge WADDR[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[5], 1.0);
   $hold(posedge WCLK, negedge WADDR[5], 1.0);
   $setup(posedge WADDR[6], posedge WCLK, 1.0);
   $setup(negedge WADDR[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[6], 1.0);
   $hold(posedge WCLK, negedge WADDR[6], 1.0);
   $setup(posedge WADDR[7], posedge WCLK, 1.0);
   $setup(negedge WADDR[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[7], 1.0);
   $hold(posedge WCLK, negedge WADDR[7], 1.0);
   $setup(posedge WADDR[8], posedge WCLK, 1.0);
   $setup(negedge WADDR[8], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[8], 1.0);
   $hold(posedge WCLK, negedge WADDR[8], 1.0);
   $setup(posedge WADDR[9], posedge WCLK, 1.0);
   $setup(negedge WADDR[9], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[9], 1.0);
   $hold(posedge WCLK, negedge WADDR[9], 1.0);
   $setup(posedge WDATA[0], posedge WCLK, 1.0);
   $setup(negedge WDATA[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[0], 1.0);
   $hold(posedge WCLK, negedge WDATA[0], 1.0);
   $setup(posedge WDATA[1], posedge WCLK, 1.0);
   $setup(negedge WDATA[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[1], 1.0);
   $hold(posedge WCLK, negedge WDATA[1], 1.0);
   $setup(posedge WDATA[2], posedge WCLK, 1.0);
   $setup(negedge WDATA[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[2], 1.0);
   $hold(posedge WCLK, negedge WDATA[2], 1.0);
   $setup(posedge WDATA[3], posedge WCLK, 1.0);
   $setup(negedge WDATA[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[3], 1.0);
   $hold(posedge WCLK, negedge WDATA[3], 1.0);
   $setup(posedge WCLKE, posedge WCLK, 1.0);
   $setup(negedge WCLKE, posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WCLKE, 1.0);
   $hold(posedge WCLK, negedge WCLKE, 1.0);
   $setup(posedge WE, posedge WCLK, 1.0);
   $setup(negedge WE, posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WE, 1.0);
   $hold(posedge WCLK, negedge WE, 1.0);
   $setup(posedge RADDR[0], posedge RCLKN, 1.0);
   $setup(negedge RADDR[0], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[0], 1.0);
   $hold(posedge RCLKN, negedge RADDR[0], 1.0);
   $setup(posedge RADDR[1], posedge RCLKN, 1.0);
   $setup(negedge RADDR[1], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[1], 1.0);
   $hold(posedge RCLKN, negedge RADDR[1], 1.0);
   $setup(posedge RADDR[2], posedge RCLKN, 1.0);
   $setup(negedge RADDR[2], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[2], 1.0);
   $hold(posedge RCLKN, negedge RADDR[2], 1.0);
   $setup(posedge RADDR[3], posedge RCLKN, 1.0);
   $setup(negedge RADDR[3], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[3], 1.0);
   $hold(posedge RCLKN, negedge RADDR[3], 1.0);
   $setup(posedge RADDR[4], posedge RCLKN, 1.0);
   $setup(negedge RADDR[4], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[4], 1.0);
   $hold(posedge RCLKN, negedge RADDR[4], 1.0);
   $setup(posedge RADDR[5], posedge RCLKN, 1.0);
   $setup(negedge RADDR[5], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[5], 1.0);
   $hold(posedge RCLKN, negedge RADDR[5], 1.0);
   $setup(posedge RADDR[6], posedge RCLKN, 1.0);
   $setup(negedge RADDR[6], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[6], 1.0);
   $hold(posedge RCLKN, negedge RADDR[6], 1.0);
   $setup(posedge RADDR[7], posedge RCLKN, 1.0);
   $setup(negedge RADDR[7], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[7], 1.0);
   $hold(posedge RCLKN, negedge RADDR[7], 1.0);
   $setup(posedge RADDR[8], posedge RCLKN, 1.0);
   $setup(negedge RADDR[8], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[8], 1.0);
   $hold(posedge RCLKN, negedge RADDR[8], 1.0);
   $setup(posedge RADDR[9], posedge RCLKN, 1.0);
   $setup(negedge RADDR[9], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[9], 1.0);
   $hold(posedge RCLKN, negedge RADDR[9], 1.0);
   $setup(posedge RCLKE, posedge RCLKN, 1.0);
   $setup(negedge RCLKE, posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RCLKE, 1.0);
   $hold(posedge RCLKN, negedge RCLKE, 1.0);
   $setup(posedge RE, posedge RCLKN, 1.0);
   $setup(negedge RE, posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RE, 1.0);
   $hold(posedge RCLKN, negedge RE, 1.0);
   $recovery(posedge RCLKN, posedge WCLK, 1.0);
   $recovery(negedge RCLKN, posedge WCLK, 1.0);
   $removal(posedge RCLKN, posedge WCLK, 1.0);
   $removal(negedge RCLKN, posedge WCLK, 1.0);
   $recovery(posedge WCLK, posedge RCLKN, 1.0);
   $recovery(negedge WCLK, posedge RCLKN, 1.0);
   $removal(posedge WCLK, posedge RCLKN, 1.0);
   $removal(negedge WCLK, posedge RCLKN, 1.0);
endspecify
`endif

endmodule //SB_RAM1024x4NR


`timescale 1ps/1ps
module SB_RAM1024x4NW (RDATA, RCLK, RCLKE, RE, RADDR, WCLKN, WCLKE, WE, WADDR, WDATA);
output [3:0] RDATA;
input RCLK;
input RCLKE;
input RE;
input [9:0] RADDR;
input WCLKN;
input WCLKE;
input WE;
input [9:0] WADDR;
input [3:0] WDATA;

parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

wire WCLK;
assign (weak0, weak1) RCLKE =1'b1 ;
assign (weak0, weak1) RE =1'b0 ;
assign (weak0, weak1) WCLKE =1'b1 ;
assign (weak0, weak1) WE =1'b0 ;
assign WCLK = ~WCLKN;

SB_RAM1024x4 sb_ram1024X4w_inst (
	.RDATA(RDATA),
	.RCLK(RCLK),
	.RCLKE(RCLKE),
	.RE(RE),
	.RADDR(RADDR),
	.WCLK(WCLK),
	.WCLKE(WCLKE),
	.WE(WE),
	.WADDR(WADDR),
	.WDATA(WDATA));

defparam sb_ram1024X4w_inst.INIT_0 = INIT_0;
defparam sb_ram1024X4w_inst.INIT_1 = INIT_1;
defparam sb_ram1024X4w_inst.INIT_2 = INIT_2;
defparam sb_ram1024X4w_inst.INIT_3 = INIT_3;
defparam sb_ram1024X4w_inst.INIT_4 = INIT_4;
defparam sb_ram1024X4w_inst.INIT_5 = INIT_5;
defparam sb_ram1024X4w_inst.INIT_6 = INIT_6;
defparam sb_ram1024X4w_inst.INIT_7 = INIT_7;
defparam sb_ram1024X4w_inst.INIT_8 = INIT_8;
defparam sb_ram1024X4w_inst.INIT_9 = INIT_9;
defparam sb_ram1024X4w_inst.INIT_A = INIT_A;
defparam sb_ram1024X4w_inst.INIT_B = INIT_B;
defparam sb_ram1024X4w_inst.INIT_C = INIT_C;
defparam sb_ram1024X4w_inst.INIT_D = INIT_D;
defparam sb_ram1024X4w_inst.INIT_E = INIT_E;
defparam sb_ram1024X4w_inst.INIT_F = INIT_F;

`ifdef TIMINGCHECK
specify
   (RCLK *> RDATA[0]) = (1.0, 1.0);
   (RCLK *> RDATA[1]) = (1.0, 1.0);
   (RCLK *> RDATA[2]) = (1.0, 1.0);
   (RCLK *> RDATA[3]) = (1.0, 1.0);
   $setup(posedge WADDR[0], posedge WCLKN, 1.0);
   $setup(negedge WADDR[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[0], 1.0);
   $hold(posedge WCLKN, negedge WADDR[0], 1.0);
   $setup(posedge WADDR[1], posedge WCLKN, 1.0);
   $setup(negedge WADDR[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[1], 1.0);
   $hold(posedge WCLKN, negedge WADDR[1], 1.0);
   $setup(posedge WADDR[2], posedge WCLKN, 1.0);
   $setup(negedge WADDR[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[2], 1.0);
   $hold(posedge WCLKN, negedge WADDR[2], 1.0);
   $setup(posedge WADDR[3], posedge WCLKN, 1.0);
   $setup(negedge WADDR[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[3], 1.0);
   $hold(posedge WCLKN, negedge WADDR[3], 1.0);
   $setup(posedge WADDR[4], posedge WCLKN, 1.0);
   $setup(negedge WADDR[4], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[4], 1.0);
   $hold(posedge WCLKN, negedge WADDR[4], 1.0);
   $setup(posedge WADDR[5], posedge WCLKN, 1.0);
   $setup(negedge WADDR[5], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[5], 1.0);
   $hold(posedge WCLKN, negedge WADDR[5], 1.0);
   $setup(posedge WADDR[6], posedge WCLKN, 1.0);
   $setup(negedge WADDR[6], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[6], 1.0);
   $hold(posedge WCLKN, negedge WADDR[6], 1.0);
   $setup(posedge WADDR[7], posedge WCLKN, 1.0);
   $setup(negedge WADDR[7], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[7], 1.0);
   $hold(posedge WCLKN, negedge WADDR[7], 1.0);
   $setup(posedge WADDR[8], posedge WCLKN, 1.0);
   $setup(negedge WADDR[8], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[8], 1.0);
   $hold(posedge WCLKN, negedge WADDR[8], 1.0);
   $setup(posedge WADDR[9], posedge WCLKN, 1.0);
   $setup(negedge WADDR[9], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[9], 1.0);
   $hold(posedge WCLKN, negedge WADDR[9], 1.0);
   $setup(posedge WDATA[0], posedge WCLKN, 1.0);
   $setup(negedge WDATA[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[0], 1.0);
   $hold(posedge WCLKN, negedge WDATA[0], 1.0);
   $setup(posedge WDATA[1], posedge WCLKN, 1.0);
   $setup(negedge WDATA[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[1], 1.0);
   $hold(posedge WCLKN, negedge WDATA[1], 1.0);
   $setup(posedge WDATA[2], posedge WCLKN, 1.0);
   $setup(negedge WDATA[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[2], 1.0);
   $hold(posedge WCLKN, negedge WDATA[2], 1.0);
   $setup(posedge WDATA[3], posedge WCLKN, 1.0);
   $setup(negedge WDATA[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[3], 1.0);
   $hold(posedge WCLKN, negedge WDATA[3], 1.0);
   $setup(posedge WCLKE, posedge WCLKN, 1.0);
   $setup(negedge WCLKE, posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WCLKE, 1.0);
   $hold(posedge WCLKN, negedge WCLKE, 1.0);
   $setup(posedge WE, posedge WCLKN, 1.0);
   $setup(negedge WE, posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WE, 1.0);
   $hold(posedge WCLKN, negedge WE, 1.0);
   $setup(posedge RADDR[0], posedge RCLK, 1.0);
   $setup(negedge RADDR[0], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[0], 1.0);
   $hold(posedge RCLK, negedge RADDR[0], 1.0);
   $setup(posedge RADDR[1], posedge RCLK, 1.0);
   $setup(negedge RADDR[1], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[1], 1.0);
   $hold(posedge RCLK, negedge RADDR[1], 1.0);
   $setup(posedge RADDR[2], posedge RCLK, 1.0);
   $setup(negedge RADDR[2], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[2], 1.0);
   $hold(posedge RCLK, negedge RADDR[2], 1.0);
   $setup(posedge RADDR[3], posedge RCLK, 1.0);
   $setup(negedge RADDR[3], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[3], 1.0);
   $hold(posedge RCLK, negedge RADDR[3], 1.0);
   $setup(posedge RADDR[4], posedge RCLK, 1.0);
   $setup(negedge RADDR[4], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[4], 1.0);
   $hold(posedge RCLK, negedge RADDR[4], 1.0);
   $setup(posedge RADDR[5], posedge RCLK, 1.0);
   $setup(negedge RADDR[5], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[5], 1.0);
   $hold(posedge RCLK, negedge RADDR[5], 1.0);
   $setup(posedge RADDR[6], posedge RCLK, 1.0);
   $setup(negedge RADDR[6], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[6], 1.0);
   $hold(posedge RCLK, negedge RADDR[6], 1.0);
   $setup(posedge RADDR[7], posedge RCLK, 1.0);
   $setup(negedge RADDR[7], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[7], 1.0);
   $hold(posedge RCLK, negedge RADDR[7], 1.0);
   $setup(posedge RADDR[8], posedge RCLK, 1.0);
   $setup(negedge RADDR[8], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[8], 1.0);
   $hold(posedge RCLK, negedge RADDR[8], 1.0);
   $setup(posedge RADDR[9], posedge RCLK, 1.0);
   $setup(negedge RADDR[9], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[9], 1.0);
   $hold(posedge RCLK, negedge RADDR[9], 1.0);
   $setup(posedge RCLKE, posedge RCLK, 1.0);
   $setup(negedge RCLKE, posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RCLKE, 1.0);
   $hold(posedge RCLK, negedge RCLKE, 1.0);
   $setup(posedge RE, posedge RCLK, 1.0);
   $setup(negedge RE, posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RE, 1.0);
   $hold(posedge RCLK, negedge RE, 1.0);
   $recovery(posedge RCLK, posedge WCLKN, 1.0);
   $recovery(negedge RCLK, posedge WCLKN, 1.0);
   $removal(posedge RCLK, posedge WCLKN, 1.0);
   $removal(negedge RCLK, posedge WCLKN, 1.0);
   $recovery(posedge WCLKN, posedge RCLK, 1.0);
   $recovery(negedge WCLKN, posedge RCLK, 1.0);
   $removal(posedge WCLKN, posedge RCLK, 1.0);
   $removal(negedge WCLKN, posedge RCLK, 1.0);

endspecify
`endif


endmodule //SB_RAM1024x4NW



`timescale 1ps/1ps
module SB_RAM1024x4NRNW (RDATA, RCLKN, RCLKE, RE, RADDR, WCLKN, WCLKE, WE, WADDR, WDATA);
output [3:0] RDATA;
input RCLKN;
input RCLKE;
input RE;
input [9:0] RADDR;
input WCLKN;
input WCLKE;
input WE;
input [9:0] WADDR;
input [3:0] WDATA;

parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

wire RCLK, WCLK;
assign (weak0, weak1) RCLKE =1'b1 ;
assign (weak0, weak1) RE =1'b0 ;
assign (weak0, weak1) WCLKE =1'b1 ;
assign (weak0, weak1) WE =1'b0 ;
assign RCLK = ~RCLKN;
assign WCLK = ~WCLKN;

SB_RAM1024x4 sb_ram1024X4rw_inst (
	.RDATA(RDATA),
	.RCLK(RCLK),
	.RCLKE(RCLKE),
	.RE(RE),
	.RADDR(RADDR),
	.WCLK(WCLK),
	.WCLKE(WCLKE),
	.WE(WE),
	.WADDR(WADDR),
	.WDATA(WDATA));

defparam sb_ram1024X4rw_inst.INIT_0 = INIT_0;
defparam sb_ram1024X4rw_inst.INIT_1 = INIT_1;
defparam sb_ram1024X4rw_inst.INIT_2 = INIT_2;
defparam sb_ram1024X4rw_inst.INIT_3 = INIT_3;
defparam sb_ram1024X4rw_inst.INIT_4 = INIT_4;
defparam sb_ram1024X4rw_inst.INIT_5 = INIT_5;
defparam sb_ram1024X4rw_inst.INIT_6 = INIT_6;
defparam sb_ram1024X4rw_inst.INIT_7 = INIT_7;
defparam sb_ram1024X4rw_inst.INIT_8 = INIT_8;
defparam sb_ram1024X4rw_inst.INIT_9 = INIT_9;
defparam sb_ram1024X4rw_inst.INIT_A = INIT_A;
defparam sb_ram1024X4rw_inst.INIT_B = INIT_B;
defparam sb_ram1024X4rw_inst.INIT_C = INIT_C;
defparam sb_ram1024X4rw_inst.INIT_D = INIT_D;
defparam sb_ram1024X4rw_inst.INIT_E = INIT_E;
defparam sb_ram1024X4rw_inst.INIT_F = INIT_F;

`ifdef TIMINGCHECK
specify
   (RCLKN *> RDATA[0]) = (1.0, 1.0);
   (RCLKN *> RDATA[1]) = (1.0, 1.0);
   (RCLKN *> RDATA[2]) = (1.0, 1.0);
   (RCLKN *> RDATA[3]) = (1.0, 1.0);
   $setup(posedge WADDR[0], posedge WCLKN, 1.0);
   $setup(negedge WADDR[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[0], 1.0);
   $hold(posedge WCLKN, negedge WADDR[0], 1.0);
   $setup(posedge WADDR[1], posedge WCLKN, 1.0);
   $setup(negedge WADDR[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[1], 1.0);
   $hold(posedge WCLKN, negedge WADDR[1], 1.0);
   $setup(posedge WADDR[2], posedge WCLKN, 1.0);
   $setup(negedge WADDR[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[2], 1.0);
   $hold(posedge WCLKN, negedge WADDR[2], 1.0);
   $setup(posedge WADDR[3], posedge WCLKN, 1.0);
   $setup(negedge WADDR[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[3], 1.0);
   $hold(posedge WCLKN, negedge WADDR[3], 1.0);
   $setup(posedge WADDR[4], posedge WCLKN, 1.0);
   $setup(negedge WADDR[4], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[4], 1.0);
   $hold(posedge WCLKN, negedge WADDR[4], 1.0);
   $setup(posedge WADDR[5], posedge WCLKN, 1.0);
   $setup(negedge WADDR[5], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[5], 1.0);
   $hold(posedge WCLKN, negedge WADDR[5], 1.0);
   $setup(posedge WADDR[6], posedge WCLKN, 1.0);
   $setup(negedge WADDR[6], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[6], 1.0);
   $hold(posedge WCLKN, negedge WADDR[6], 1.0);
   $setup(posedge WADDR[7], posedge WCLKN, 1.0);
   $setup(negedge WADDR[7], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[7], 1.0);
   $hold(posedge WCLKN, negedge WADDR[7], 1.0);
   $setup(posedge WADDR[8], posedge WCLKN, 1.0);
   $setup(negedge WADDR[8], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[8], 1.0);
   $hold(posedge WCLKN, negedge WADDR[8], 1.0);
   $setup(posedge WADDR[9], posedge WCLKN, 1.0);
   $setup(negedge WADDR[9], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[9], 1.0);
   $hold(posedge WCLKN, negedge WADDR[9], 1.0);
   $setup(posedge WDATA[0], posedge WCLKN, 1.0);
   $setup(negedge WDATA[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[0], 1.0);
   $hold(posedge WCLKN, negedge WDATA[0], 1.0);
   $setup(posedge WDATA[1], posedge WCLKN, 1.0);
   $setup(negedge WDATA[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[1], 1.0);
   $hold(posedge WCLKN, negedge WDATA[1], 1.0);
   $setup(posedge WDATA[2], posedge WCLKN, 1.0);
   $setup(negedge WDATA[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[2], 1.0);
   $hold(posedge WCLKN, negedge WDATA[2], 1.0);
   $setup(posedge WDATA[3], posedge WCLKN, 1.0);
   $setup(negedge WDATA[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[3], 1.0);
   $hold(posedge WCLKN, negedge WDATA[3], 1.0);
   $setup(posedge WCLKE, posedge WCLKN, 1.0);
   $setup(negedge WCLKE, posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WCLKE, 1.0);
   $hold(posedge WCLKN, negedge WCLKE, 1.0);
   $setup(posedge WE, posedge WCLKN, 1.0);
   $setup(negedge WE, posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WE, 1.0);
   $hold(posedge WCLKN, negedge WE, 1.0);
   $setup(posedge RADDR[0], posedge RCLKN, 1.0);
   $setup(negedge RADDR[0], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[0], 1.0);
   $hold(posedge RCLKN, negedge RADDR[0], 1.0);
   $setup(posedge RADDR[1], posedge RCLKN, 1.0);
   $setup(negedge RADDR[1], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[1], 1.0);
   $hold(posedge RCLKN, negedge RADDR[1], 1.0);
   $setup(posedge RADDR[2], posedge RCLKN, 1.0);
   $setup(negedge RADDR[2], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[2], 1.0);
   $hold(posedge RCLKN, negedge RADDR[2], 1.0);
   $setup(posedge RADDR[3], posedge RCLKN, 1.0);
   $setup(negedge RADDR[3], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[3], 1.0);
   $hold(posedge RCLKN, negedge RADDR[3], 1.0);
   $setup(posedge RADDR[4], posedge RCLKN, 1.0);
   $setup(negedge RADDR[4], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[4], 1.0);
   $hold(posedge RCLKN, negedge RADDR[4], 1.0);
   $setup(posedge RADDR[5], posedge RCLKN, 1.0);
   $setup(negedge RADDR[5], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[5], 1.0);
   $hold(posedge RCLKN, negedge RADDR[5], 1.0);
   $setup(posedge RADDR[6], posedge RCLKN, 1.0);
   $setup(negedge RADDR[6], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[6], 1.0);
   $hold(posedge RCLKN, negedge RADDR[6], 1.0);
   $setup(posedge RADDR[7], posedge RCLKN, 1.0);
   $setup(negedge RADDR[7], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[7], 1.0);
   $hold(posedge RCLKN, negedge RADDR[7], 1.0);
   $setup(posedge RADDR[8], posedge RCLKN, 1.0);
   $setup(negedge RADDR[8], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[8], 1.0);
   $hold(posedge RCLKN, negedge RADDR[8], 1.0);
   $setup(posedge RADDR[9], posedge RCLKN, 1.0);
   $setup(negedge RADDR[9], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[9], 1.0);
   $hold(posedge RCLKN, negedge RADDR[9], 1.0);
   $setup(posedge RCLKE, posedge RCLKN, 1.0);
   $setup(negedge RCLKE, posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RCLKE, 1.0);
   $hold(posedge RCLKN, negedge RCLKE, 1.0);
   $setup(posedge RE, posedge RCLKN, 1.0);
   $setup(negedge RE, posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RE, 1.0);
   $hold(posedge RCLKN, negedge RE, 1.0);
   $recovery(posedge RCLKN, posedge WCLKN, 1.0);
   $recovery(negedge RCLKN, posedge WCLKN, 1.0);
   $removal(posedge RCLKN, posedge WCLKN, 1.0);
   $removal(negedge RCLKN, posedge WCLKN, 1.0);
   $recovery(posedge WCLKN, posedge RCLKN, 1.0);
   $recovery(negedge WCLKN, posedge RCLKN, 1.0);
   $removal(posedge WCLKN, posedge RCLKN, 1.0);
   $removal(negedge WCLKN, posedge RCLKN, 1.0);

endspecify
`endif
endmodule //SB_RAM1024x4NRNW



`timescale 1ps/1ps
module SB_RAM2048x2 (RDATA, RCLK, RCLKE, RE, RADDR, WCLK, WCLKE, WE, WADDR, WDATA);
output [1:0] RDATA;
input RCLK;
input RCLKE;
input RE;
input [10:0] RADDR;
input WCLK;
input WCLKE;
input WE;
input [10:0] WADDR;
input [1:0] WDATA;

parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

// local Parameters
localparam			CLOCK_PERIOD = 200;	//
localparam 			DELAY	= (CLOCK_PERIOD/10);		// Clock-to-output delay. Zero
							// time delays can be confusing
							// and sometimes cause problems.
localparam 			BUS_WIDTH = 2;		// Width of RAM (number of bits)

localparam 			ADDRESS_BUS_SIZE = 11;	// Number of bits required to
							// represent the RAM address

localparam   ADDRESSABLE_SPACE  = 2**ADDRESS_BUS_SIZE;	// Decimal address range [2^Size:0]


// SIGNAL DECLARATIONS
wire			   	WCLK_g, RCLK_g;
reg 				WCLKE_sync, RCLKE_sync; 
assign (weak0, weak1) RCLKE =1'b1 ;
assign (weak0, weak1) RE =1'b0 ;
assign (weak0, weak1) WCLKE =1'b1 ;
assign (weak0, weak1) WE =1'b0 ;
reg	Memory	[BUS_WIDTH*ADDRESSABLE_SPACE-1:0];
// 
event Read_e, Write_e;

//////////////////// Collision detect begins here ///////////////////////////////
localparam 	TRUE = 1'b1;
localparam	FALSE = 1'b0;
reg 		Time_Collision_Detected = 1'b0;
wire		Address_Collision_Detected;

event Collision_e;

time COLLISION_TIME_WINDOW = (CLOCK_PERIOD/8); // This is an arbitray value, but is better than using an absolute 
						    // value, because the actual time window depends on the actual silicon 
						    // implementation. Thus the test is indicative of an Error and not
						    // guaranteed to be an error. Even so this is usefull.
time time_WCLK_RCLK, time_WCLK, time_RCLK;


//function reg Check_Timed_Window_Violation;
function	Check_Timed_Window_Violation;	//	by Jeffrey
input T1, T2, Minimum_Time_Window;
time T1, T2;
time Minimum_Time_Window;
time Difference;	
	begin
		Difference = (T1 - T2);
		if (Difference < 0) Difference = -Difference;
		Check_Timed_Window_Violation = (Difference < Minimum_Time_Window);
	end
endfunction


initial begin
       time_WCLK = CLOCK_PERIOD;	// Arbitrary initialisation value, ensure no window collison error on first clock edge.
       time_RCLK = (CLOCK_PERIOD*8);	// Arbitrary initialisation difference value, ensure no collision error on first clock edge.					
end

integer	i,j;


initial	//	initialize ram_4k by parameter, section by section
begin
	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[BUS_WIDTH*i+j]	=	INIT_0[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*1+BUS_WIDTH*i+j]	=	INIT_1[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*2+BUS_WIDTH*i+j]	=	INIT_2[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*3+BUS_WIDTH*i+j]	=	INIT_3[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*4+BUS_WIDTH*i+j]	=	INIT_4[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*5+BUS_WIDTH*i+j]	=	INIT_5[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*6+BUS_WIDTH*i+j]	=	INIT_6[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*7+BUS_WIDTH*i+j]	=	INIT_7[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*8+BUS_WIDTH*i+j]	=	INIT_8[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*9+BUS_WIDTH*i+j]	=	INIT_9[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*10+BUS_WIDTH*i+j]	=	INIT_A[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*11+BUS_WIDTH*i+j]	=	INIT_B[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*12+BUS_WIDTH*i+j]	=	INIT_C[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*13+BUS_WIDTH*i+j]	=	INIT_D[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*14+BUS_WIDTH*i+j]	=	INIT_E[BUS_WIDTH*i+j];
	end

	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
			Memory[256*15+BUS_WIDTH*i+j]	=	INIT_F[BUS_WIDTH*i+j];
	end

end

assign Address_Collision_Detected = ((RE & WE & WCLKE & RCLKE)&(WADDR == RADDR)); 

always @(WCLK or WCLKE) 
begin 
	if(~WCLK)
	WCLKE_sync = WCLKE;   	
end 

always @(RCLK or RCLKE) 
begin 
	if (~RCLK)
	RCLKE_sync = RCLKE; 	
end 

assign WCLK_g = WCLK & WCLKE_sync;
assign RCLK_g = RCLK & RCLKE_sync;

always @(posedge WCLK_g) begin
	time_WCLK = $time;
end

always @(posedge RCLK_g) begin
    	time_RCLK = $time;
end
integer	SB_RAM2048X2_RDATA_log_file;					//.....................
initial	SB_RAM2048X2_RDATA_log_file=("SB_RAM2048X2_RDATA_log_file.txt");	//.....................
always @(posedge WCLK_g) begin

	Time_Collision_Detected = Check_Timed_Window_Violation(time_WCLK,time_RCLK,COLLISION_TIME_WINDOW);
        if (Time_Collision_Detected & Address_Collision_Detected)begin
        	$display("Warning: Write-Read collision detected, Data read value is X\n");
 		$display("WCLK Time: %.3f   RCLK Time:%.3f  ",time_WCLK, time_RCLK,"WADDR: %d   RADDR:%d\n",WADDR, RADDR); 
 		$fdisplay(SB_RAM2048X2_RDATA_log_file,"Warning: Write-Read collision detected, Data read value is X\n");
		$fdisplay(SB_RAM2048X2_RDATA_log_file,"WCLK Time: %.3f   RCLK Time:%.3f  ",time_WCLK, time_RCLK, "WADDR: %d   RADDR:%d\n",WADDR, RADDR); 	
 		-> Collision_e;
	end
end




//	code modify for universal verilog compiler

always @ (posedge WCLK_g)
begin
	if	(WE)
	begin
		-> Write_e;
		for	(i=0;i<=BUS_WIDTH-1; i=i+1)
		begin
			Memory[WADDR*BUS_WIDTH+i]	<=	WDATA[i];
		end
	end
end

//reg	[1:0]	RDATA = 0;
reg	[1:0]	RDATA = 0;

initial
begin
   RDATA = $random;
end

// Look at the rising edge of the clock

always @ (posedge RCLK_g)
begin
	if	(RE)
	begin
		-> Read_e;
		if	(Time_Collision_Detected & Address_Collision_Detected) 
			RDATA <= 2'hX;
		else
			for	(i=0;i<=BUS_WIDTH-1;i=i+1)
				RDATA[i]	<= Memory[RADDR*BUS_WIDTH+i];
	end
end

`ifdef TIMINGCHECK
specify
   (RCLK *> RDATA[0]) = (1.0, 1.0);
   (RCLK *> RDATA[1]) = (1.0, 1.0);
   $setup(posedge WADDR[0], posedge WCLK, 1.0);
   $setup(negedge WADDR[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[0], 1.0);
   $hold(posedge WCLK, negedge WADDR[0], 1.0);
   $setup(posedge WADDR[1], posedge WCLK, 1.0);
   $setup(negedge WADDR[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[1], 1.0);
   $hold(posedge WCLK, negedge WADDR[1], 1.0);
   $setup(posedge WADDR[2], posedge WCLK, 1.0);
   $setup(negedge WADDR[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[2], 1.0);
   $hold(posedge WCLK, negedge WADDR[2], 1.0);
   $setup(posedge WADDR[3], posedge WCLK, 1.0);
   $setup(negedge WADDR[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[3], 1.0);
   $hold(posedge WCLK, negedge WADDR[3], 1.0);
   $setup(posedge WADDR[4], posedge WCLK, 1.0);
   $setup(negedge WADDR[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[4], 1.0);
   $hold(posedge WCLK, negedge WADDR[4], 1.0);
   $setup(posedge WADDR[5], posedge WCLK, 1.0);
   $setup(negedge WADDR[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[5], 1.0);
   $hold(posedge WCLK, negedge WADDR[5], 1.0);
   $setup(posedge WADDR[6], posedge WCLK, 1.0);
   $setup(negedge WADDR[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[6], 1.0);
   $hold(posedge WCLK, negedge WADDR[6], 1.0);
   $setup(posedge WADDR[7], posedge WCLK, 1.0);
   $setup(negedge WADDR[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[7], 1.0);
   $hold(posedge WCLK, negedge WADDR[7], 1.0);
   $setup(posedge WADDR[8], posedge WCLK, 1.0);
   $setup(negedge WADDR[8], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[8], 1.0);
   $hold(posedge WCLK, negedge WADDR[8], 1.0);
   $setup(posedge WADDR[9], posedge WCLK, 1.0);
   $setup(negedge WADDR[9], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[9], 1.0);
   $hold(posedge WCLK, negedge WADDR[9], 1.0);
   $setup(posedge WADDR[10], posedge WCLK, 1.0);
   $setup(negedge WADDR[10], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[10], 1.0);
   $hold(posedge WCLK, negedge WADDR[10], 1.0);
   $setup(posedge WDATA[0], posedge WCLK, 1.0);
   $setup(negedge WDATA[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[0], 1.0);
   $hold(posedge WCLK, negedge WDATA[0], 1.0);
   $setup(posedge WDATA[1], posedge WCLK, 1.0);
   $setup(negedge WDATA[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[1], 1.0);
   $hold(posedge WCLK, negedge WDATA[1], 1.0);
   $setup(posedge WCLKE, posedge WCLK, 1.0);
   $setup(negedge WCLKE, posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WCLKE, 1.0);
   $hold(posedge WCLK, negedge WCLKE, 1.0);
   $setup(posedge WE, posedge WCLK, 1.0);
   $setup(negedge WE, posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WE, 1.0);
   $hold(posedge WCLK, negedge WE, 1.0);
   $setup(posedge RADDR[0], posedge RCLK, 1.0);
   $setup(negedge RADDR[0], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[0], 1.0);
   $hold(posedge RCLK, negedge RADDR[0], 1.0);
   $setup(posedge RADDR[1], posedge RCLK, 1.0);
   $setup(negedge RADDR[1], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[1], 1.0);
   $hold(posedge RCLK, negedge RADDR[1], 1.0);
   $setup(posedge RADDR[2], posedge RCLK, 1.0);
   $setup(negedge RADDR[2], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[2], 1.0);
   $hold(posedge RCLK, negedge RADDR[2], 1.0);
   $setup(posedge RADDR[3], posedge RCLK, 1.0);
   $setup(negedge RADDR[3], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[3], 1.0);
   $hold(posedge RCLK, negedge RADDR[3], 1.0);
   $setup(posedge RADDR[4], posedge RCLK, 1.0);
   $setup(negedge RADDR[4], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[4], 1.0);
   $hold(posedge RCLK, negedge RADDR[4], 1.0);
   $setup(posedge RADDR[5], posedge RCLK, 1.0);
   $setup(negedge RADDR[5], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[5], 1.0);
   $hold(posedge RCLK, negedge RADDR[5], 1.0);
   $setup(posedge RADDR[6], posedge RCLK, 1.0);
   $setup(negedge RADDR[6], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[6], 1.0);
   $hold(posedge RCLK, negedge RADDR[6], 1.0);
   $setup(posedge RADDR[7], posedge RCLK, 1.0);
   $setup(negedge RADDR[7], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[7], 1.0);
   $hold(posedge RCLK, negedge RADDR[7], 1.0);
   $setup(posedge RADDR[8], posedge RCLK, 1.0);
   $setup(negedge RADDR[8], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[8], 1.0);
   $hold(posedge RCLK, negedge RADDR[8], 1.0);
   $setup(posedge RADDR[9], posedge RCLK, 1.0);
   $setup(negedge RADDR[9], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[9], 1.0);
   $hold(posedge RCLK, negedge RADDR[9], 1.0);
   $setup(posedge RADDR[10], posedge RCLK, 1.0);
   $setup(negedge RADDR[10], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[10], 1.0);
   $hold(posedge RCLK, negedge RADDR[10], 1.0);
   $setup(posedge RCLKE, posedge RCLK, 1.0);
   $setup(negedge RCLKE, posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RCLKE, 1.0);
   $hold(posedge RCLK, negedge RCLKE, 1.0);
   $setup(posedge RE, posedge RCLK, 1.0);
   $setup(negedge RE, posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RE, 1.0);
   $hold(posedge RCLK, negedge RE, 1.0);

endspecify
`endif
endmodule //SB_RAM2048x2


`timescale 1ps/1ps
module SB_RAM2048x2NR (RDATA, RCLKN, RCLKE, RE, RADDR, WCLK, WCLKE, WE, WADDR, WDATA);
output [1:0] RDATA;
input RCLKN;
input RCLKE;
input RE;
input [10:0] RADDR;
input WCLK;
input WCLKE;
input WE;
input [10:0] WADDR;
input [1:0] WDATA;

parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

wire RCLK;
assign (weak0, weak1) RCLKE =1'b1 ;
assign (weak0, weak1) RE =1'b0 ;
assign (weak0, weak1) WCLKE =1'b1 ;
assign (weak0, weak1) WE =1'b0 ;
assign RCLK = ~RCLKN;

SB_RAM2048x2 sb_ram2048X2r_inst (
	.RDATA(RDATA),
	.RCLK(RCLK),
	.RCLKE(RCLKE),
	.RE(RE),
	.RADDR(RADDR),
	.WCLK(WCLK),
	.WCLKE(WCLKE),
	.WE(WE),
	.WADDR(WADDR),
	.WDATA(WDATA));

defparam sb_ram2048X2r_inst.INIT_0 = INIT_0;
defparam sb_ram2048X2r_inst.INIT_1 = INIT_1;
defparam sb_ram2048X2r_inst.INIT_2 = INIT_2;
defparam sb_ram2048X2r_inst.INIT_3 = INIT_3;
defparam sb_ram2048X2r_inst.INIT_4 = INIT_4;
defparam sb_ram2048X2r_inst.INIT_5 = INIT_5;
defparam sb_ram2048X2r_inst.INIT_6 = INIT_6;
defparam sb_ram2048X2r_inst.INIT_7 = INIT_7;
defparam sb_ram2048X2r_inst.INIT_8 = INIT_8;
defparam sb_ram2048X2r_inst.INIT_9 = INIT_9;
defparam sb_ram2048X2r_inst.INIT_A = INIT_A;
defparam sb_ram2048X2r_inst.INIT_B = INIT_B;
defparam sb_ram2048X2r_inst.INIT_C = INIT_C;
defparam sb_ram2048X2r_inst.INIT_D = INIT_D;
defparam sb_ram2048X2r_inst.INIT_E = INIT_E;
defparam sb_ram2048X2r_inst.INIT_F = INIT_F;

`ifdef TIMINGCHECK
specify
   (RCLKN *> RDATA[0]) = (1.0, 1.0);
   (RCLKN *> RDATA[1]) = (1.0, 1.0);
   $setup(posedge WADDR[0], posedge WCLK, 1.0);
   $setup(negedge WADDR[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[0], 1.0);
   $hold(posedge WCLK, negedge WADDR[0], 1.0);
   $setup(posedge WADDR[1], posedge WCLK, 1.0);
   $setup(negedge WADDR[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[1], 1.0);
   $hold(posedge WCLK, negedge WADDR[1], 1.0);
   $setup(posedge WADDR[2], posedge WCLK, 1.0);
   $setup(negedge WADDR[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[2], 1.0);
   $hold(posedge WCLK, negedge WADDR[2], 1.0);
   $setup(posedge WADDR[3], posedge WCLK, 1.0);
   $setup(negedge WADDR[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[3], 1.0);
   $hold(posedge WCLK, negedge WADDR[3], 1.0);
   $setup(posedge WADDR[4], posedge WCLK, 1.0);
   $setup(negedge WADDR[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[4], 1.0);
   $hold(posedge WCLK, negedge WADDR[4], 1.0);
   $setup(posedge WADDR[5], posedge WCLK, 1.0);
   $setup(negedge WADDR[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[5], 1.0);
   $hold(posedge WCLK, negedge WADDR[5], 1.0);
   $setup(posedge WADDR[6], posedge WCLK, 1.0);
   $setup(negedge WADDR[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[6], 1.0);
   $hold(posedge WCLK, negedge WADDR[6], 1.0);
   $setup(posedge WADDR[7], posedge WCLK, 1.0);
   $setup(negedge WADDR[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[7], 1.0);
   $hold(posedge WCLK, negedge WADDR[7], 1.0);
   $setup(posedge WADDR[8], posedge WCLK, 1.0);
   $setup(negedge WADDR[8], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[8], 1.0);
   $hold(posedge WCLK, negedge WADDR[8], 1.0);
   $setup(posedge WADDR[9], posedge WCLK, 1.0);
   $setup(negedge WADDR[9], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[9], 1.0);
   $hold(posedge WCLK, negedge WADDR[9], 1.0);
   $setup(posedge WADDR[10], posedge WCLK, 1.0);
   $setup(negedge WADDR[10], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[10], 1.0);
   $hold(posedge WCLK, negedge WADDR[10], 1.0);
   $setup(posedge WDATA[0], posedge WCLK, 1.0);
   $setup(negedge WDATA[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[0], 1.0);
   $hold(posedge WCLK, negedge WDATA[0], 1.0);
   $setup(posedge WDATA[1], posedge WCLK, 1.0);
   $setup(negedge WDATA[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[1], 1.0);
   $hold(posedge WCLK, negedge WDATA[1], 1.0);
   $setup(posedge WCLKE, posedge WCLK, 1.0);
   $setup(negedge WCLKE, posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WCLKE, 1.0);
   $hold(posedge WCLK, negedge WCLKE, 1.0);
   $setup(posedge WE, posedge WCLK, 1.0);
   $setup(negedge WE, posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WE, 1.0);
   $hold(posedge WCLK, negedge WE, 1.0);
   $setup(posedge RADDR[0], posedge RCLKN, 1.0);
   $setup(negedge RADDR[0], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[0], 1.0);
   $hold(posedge RCLKN, negedge RADDR[0], 1.0);
   $setup(posedge RADDR[1], posedge RCLKN, 1.0);
   $setup(negedge RADDR[1], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[1], 1.0);
   $hold(posedge RCLKN, negedge RADDR[1], 1.0);
   $setup(posedge RADDR[2], posedge RCLKN, 1.0);
   $setup(negedge RADDR[2], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[2], 1.0);
   $hold(posedge RCLKN, negedge RADDR[2], 1.0);
   $setup(posedge RADDR[3], posedge RCLKN, 1.0);
   $setup(negedge RADDR[3], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[3], 1.0);
   $hold(posedge RCLKN, negedge RADDR[3], 1.0);
   $setup(posedge RADDR[4], posedge RCLKN, 1.0);
   $setup(negedge RADDR[4], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[4], 1.0);
   $hold(posedge RCLKN, negedge RADDR[4], 1.0);
   $setup(posedge RADDR[5], posedge RCLKN, 1.0);
   $setup(negedge RADDR[5], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[5], 1.0);
   $hold(posedge RCLKN, negedge RADDR[5], 1.0);
   $setup(posedge RADDR[6], posedge RCLKN, 1.0);
   $setup(negedge RADDR[6], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[6], 1.0);
   $hold(posedge RCLKN, negedge RADDR[6], 1.0);
   $setup(posedge RADDR[7], posedge RCLKN, 1.0);
   $setup(negedge RADDR[7], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[7], 1.0);
   $hold(posedge RCLKN, negedge RADDR[7], 1.0);
   $setup(posedge RADDR[8], posedge RCLKN, 1.0);
   $setup(negedge RADDR[8], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[8], 1.0);
   $hold(posedge RCLKN, negedge RADDR[8], 1.0);
   $setup(posedge RADDR[9], posedge RCLKN, 1.0);
   $setup(negedge RADDR[9], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[9], 1.0);
   $hold(posedge RCLKN, negedge RADDR[9], 1.0);
   $setup(posedge RADDR[10], posedge RCLKN, 1.0);
   $setup(negedge RADDR[10], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[10], 1.0);
   $hold(posedge RCLKN, negedge RADDR[10], 1.0);
   $setup(posedge RCLKE, posedge RCLKN, 1.0);
   $setup(negedge RCLKE, posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RCLKE, 1.0);
   $hold(posedge RCLKN, negedge RCLKE, 1.0);
   $setup(posedge RE, posedge RCLKN, 1.0);
   $setup(negedge RE, posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RE, 1.0);
   $hold(posedge RCLKN, negedge RE, 1.0);
   $recovery(posedge RCLKN, posedge WCLK, 1.0);
   $recovery(negedge RCLKN, posedge WCLK, 1.0);
   $removal(posedge RCLKN, posedge WCLK, 1.0);
   $removal(negedge RCLKN, posedge WCLK, 1.0);
   $recovery(posedge WCLK, posedge RCLKN, 1.0);
   $recovery(negedge WCLK, posedge RCLKN, 1.0);
   $removal(posedge WCLK, posedge RCLKN, 1.0);
   $removal(negedge WCLK, posedge RCLKN, 1.0);
endspecify
`endif

endmodule //SB_RAM2048x2NR



`timescale 1ps/1ps
module SB_RAM2048x2NW (RDATA, RCLK, RCLKE, RE, RADDR, WCLKN, WCLKE, WE, WADDR, WDATA);
output [1:0] RDATA;
input RCLK;
input RCLKE;
input RE;
input [10:0] RADDR;
input WCLKN;
input WCLKE;
input WE;
input [10:0] WADDR;
input [1:0] WDATA;

parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;


wire WCLK;
assign (weak0, weak1) RCLKE =1'b1 ;
assign (weak0, weak1) RE =1'b0 ;
assign (weak0, weak1) WCLKE =1'b1 ;
assign (weak0, weak1) WE =1'b0 ;
assign WCLK = ~WCLKN;

SB_RAM2048x2 sb_ram2048X2w_inst (
	.RDATA(RDATA),
	.RCLK(RCLK),
	.RCLKE(RCLKE),
	.RE(RE),
	.RADDR(RADDR),
	.WCLK(WCLK),
	.WCLKE(WCLKE),
	.WE(WE),
	.WADDR(WADDR),
	.WDATA(WDATA));

defparam sb_ram2048X2w_inst.INIT_0 = INIT_0;
defparam sb_ram2048X2w_inst.INIT_1 = INIT_1;
defparam sb_ram2048X2w_inst.INIT_2 = INIT_2;
defparam sb_ram2048X2w_inst.INIT_3 = INIT_3;
defparam sb_ram2048X2w_inst.INIT_4 = INIT_4;
defparam sb_ram2048X2w_inst.INIT_5 = INIT_5;
defparam sb_ram2048X2w_inst.INIT_6 = INIT_6;
defparam sb_ram2048X2w_inst.INIT_7 = INIT_7;
defparam sb_ram2048X2w_inst.INIT_8 = INIT_8;
defparam sb_ram2048X2w_inst.INIT_9 = INIT_9;
defparam sb_ram2048X2w_inst.INIT_A = INIT_A;
defparam sb_ram2048X2w_inst.INIT_B = INIT_B;
defparam sb_ram2048X2w_inst.INIT_C = INIT_C;
defparam sb_ram2048X2w_inst.INIT_D = INIT_D;
defparam sb_ram2048X2w_inst.INIT_E = INIT_E;
defparam sb_ram2048X2w_inst.INIT_F = INIT_F;

`ifdef TIMINGCHECK
specify
   (RCLK *> RDATA[0]) = (1.0, 1.0);
   (RCLK *> RDATA[1]) = (1.0, 1.0);
   $setup(posedge WADDR[0], posedge WCLKN, 1.0);
   $setup(negedge WADDR[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[0], 1.0);
   $hold(posedge WCLKN, negedge WADDR[0], 1.0);
   $setup(posedge WADDR[1], posedge WCLKN, 1.0);
   $setup(negedge WADDR[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[1], 1.0);
   $hold(posedge WCLKN, negedge WADDR[1], 1.0);
   $setup(posedge WADDR[2], posedge WCLKN, 1.0);
   $setup(negedge WADDR[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[2], 1.0);
   $hold(posedge WCLKN, negedge WADDR[2], 1.0);
   $setup(posedge WADDR[3], posedge WCLKN, 1.0);
   $setup(negedge WADDR[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[3], 1.0);
   $hold(posedge WCLKN, negedge WADDR[3], 1.0);
   $setup(posedge WADDR[4], posedge WCLKN, 1.0);
   $setup(negedge WADDR[4], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[4], 1.0);
   $hold(posedge WCLKN, negedge WADDR[4], 1.0);
   $setup(posedge WADDR[5], posedge WCLKN, 1.0);
   $setup(negedge WADDR[5], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[5], 1.0);
   $hold(posedge WCLKN, negedge WADDR[5], 1.0);
   $setup(posedge WADDR[6], posedge WCLKN, 1.0);
   $setup(negedge WADDR[6], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[6], 1.0);
   $hold(posedge WCLKN, negedge WADDR[6], 1.0);
   $setup(posedge WADDR[7], posedge WCLKN, 1.0);
   $setup(negedge WADDR[7], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[7], 1.0);
   $hold(posedge WCLKN, negedge WADDR[7], 1.0);
   $setup(posedge WADDR[8], posedge WCLKN, 1.0);
   $setup(negedge WADDR[8], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[8], 1.0);
   $hold(posedge WCLKN, negedge WADDR[8], 1.0);
   $setup(posedge WADDR[9], posedge WCLKN, 1.0);
   $setup(negedge WADDR[9], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[9], 1.0);
   $hold(posedge WCLKN, negedge WADDR[9], 1.0);
   $setup(posedge WADDR[10], posedge WCLKN, 1.0);
   $setup(negedge WADDR[10], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[10], 1.0);
   $hold(posedge WCLKN, negedge WADDR[10], 1.0);
   $setup(posedge WDATA[0], posedge WCLKN, 1.0);
   $setup(negedge WDATA[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[0], 1.0);
   $hold(posedge WCLKN, negedge WDATA[0], 1.0);
   $setup(posedge WDATA[1], posedge WCLKN, 1.0);
   $setup(negedge WDATA[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[1], 1.0);
   $hold(posedge WCLKN, negedge WDATA[1], 1.0);
   $setup(posedge WCLKE, posedge WCLKN, 1.0);
   $setup(negedge WCLKE, posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WCLKE, 1.0);
   $hold(posedge WCLKN, negedge WCLKE, 1.0);
   $setup(posedge WE, posedge WCLKN, 1.0);
   $setup(negedge WE, posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WE, 1.0);
   $hold(posedge WCLKN, negedge WE, 1.0);
   $setup(posedge RADDR[0], posedge RCLK, 1.0);
   $setup(negedge RADDR[0], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[0], 1.0);
   $hold(posedge RCLK, negedge RADDR[0], 1.0);
   $setup(posedge RADDR[1], posedge RCLK, 1.0);
   $setup(negedge RADDR[1], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[1], 1.0);
   $hold(posedge RCLK, negedge RADDR[1], 1.0);
   $setup(posedge RADDR[2], posedge RCLK, 1.0);
   $setup(negedge RADDR[2], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[2], 1.0);
   $hold(posedge RCLK, negedge RADDR[2], 1.0);
   $setup(posedge RADDR[3], posedge RCLK, 1.0);
   $setup(negedge RADDR[3], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[3], 1.0);
   $hold(posedge RCLK, negedge RADDR[3], 1.0);
   $setup(posedge RADDR[4], posedge RCLK, 1.0);
   $setup(negedge RADDR[4], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[4], 1.0);
   $hold(posedge RCLK, negedge RADDR[4], 1.0);
   $setup(posedge RADDR[5], posedge RCLK, 1.0);
   $setup(negedge RADDR[5], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[5], 1.0);
   $hold(posedge RCLK, negedge RADDR[5], 1.0);
   $setup(posedge RADDR[6], posedge RCLK, 1.0);
   $setup(negedge RADDR[6], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[6], 1.0);
   $hold(posedge RCLK, negedge RADDR[6], 1.0);
   $setup(posedge RADDR[7], posedge RCLK, 1.0);
   $setup(negedge RADDR[7], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[7], 1.0);
   $hold(posedge RCLK, negedge RADDR[7], 1.0);
   $setup(posedge RADDR[8], posedge RCLK, 1.0);
   $setup(negedge RADDR[8], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[8], 1.0);
   $hold(posedge RCLK, negedge RADDR[8], 1.0);
   $setup(posedge RADDR[9], posedge RCLK, 1.0);
   $setup(negedge RADDR[9], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[9], 1.0);
   $hold(posedge RCLK, negedge RADDR[9], 1.0);
   $setup(posedge RADDR[9], posedge RCLK, 1.0);
   $setup(negedge RADDR[9], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[9], 1.0);
   $hold(posedge RCLK, negedge RADDR[9], 1.0);
   $setup(posedge RCLKE, posedge RCLK, 1.0);
   $setup(negedge RCLKE, posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RCLKE, 1.0);
   $hold(posedge RCLK, negedge RCLKE, 1.0);
   $setup(posedge RE, posedge RCLK, 1.0);
   $setup(negedge RE, posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RE, 1.0);
   $hold(posedge RCLK, negedge RE, 1.0);
   $recovery(posedge RCLK, posedge WCLKN, 1.0);
   $recovery(negedge RCLK, posedge WCLKN, 1.0);
   $removal(posedge RCLK, posedge WCLKN, 1.0);
   $removal(negedge RCLK, posedge WCLKN, 1.0);
   $recovery(posedge WCLKN, posedge RCLK, 1.0);
   $recovery(negedge WCLKN, posedge RCLK, 1.0);
   $removal(posedge WCLKN, posedge RCLK, 1.0);
   $removal(negedge WCLKN, posedge RCLK, 1.0);

endspecify
`endif
endmodule //SB_RAM2048x2NW



`timescale 1ps/1ps
module SB_RAM2048x2NRNW (RDATA, RCLKN, RCLKE, RE, RADDR, WCLKN, WCLKE, WE, WADDR, WDATA);
output [1:0] RDATA;
input RCLKN;
input RCLKE;
input RE;
input [10:0] RADDR;
input WCLKN;
input WCLKE;
input WE;
input [10:0] WADDR;
input [1:0] WDATA;

parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

wire RCLK, WCLK;
assign (weak0, weak1) RCLKE =1'b1 ;
assign (weak0, weak1) RE =1'b0 ;
assign (weak0, weak1) WCLKE =1'b1 ;
assign (weak0, weak1) WE =1'b0 ;
assign RCLK = ~RCLKN;
assign WCLK = ~WCLKN;

SB_RAM2048x2 sb_ram2048X2rw_inst (
	.RDATA(RDATA),
	.RCLK(RCLK),
	.RCLKE(RCLKE),
	.RE(RE),
	.RADDR(RADDR),
	.WCLK(WCLK),
	.WCLKE(WCLKE),
	.WE(WE),
	.WADDR(WADDR),
	.WDATA(WDATA));

defparam sb_ram2048X2rw_inst.INIT_0 = INIT_0;
defparam sb_ram2048X2rw_inst.INIT_1 = INIT_1;
defparam sb_ram2048X2rw_inst.INIT_2 = INIT_2;
defparam sb_ram2048X2rw_inst.INIT_3 = INIT_3;
defparam sb_ram2048X2rw_inst.INIT_4 = INIT_4;
defparam sb_ram2048X2rw_inst.INIT_5 = INIT_5;
defparam sb_ram2048X2rw_inst.INIT_6 = INIT_6;
defparam sb_ram2048X2rw_inst.INIT_7 = INIT_7;
defparam sb_ram2048X2rw_inst.INIT_8 = INIT_8;
defparam sb_ram2048X2rw_inst.INIT_9 = INIT_9;
defparam sb_ram2048X2rw_inst.INIT_A = INIT_A;
defparam sb_ram2048X2rw_inst.INIT_B = INIT_B;
defparam sb_ram2048X2rw_inst.INIT_C = INIT_C;
defparam sb_ram2048X2rw_inst.INIT_D = INIT_D;
defparam sb_ram2048X2rw_inst.INIT_E = INIT_E;
defparam sb_ram2048X2rw_inst.INIT_F = INIT_F;

`ifdef TIMINGCHECK
specify
   (RCLKN *> RDATA[0]) = (1.0, 1.0);
   (RCLKN *> RDATA[1]) = (1.0, 1.0);
   $setup(posedge WADDR[0], posedge WCLKN, 1.0);
   $setup(negedge WADDR[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[0], 1.0);
   $hold(posedge WCLKN, negedge WADDR[0], 1.0);
   $setup(posedge WADDR[1], posedge WCLKN, 1.0);
   $setup(negedge WADDR[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[1], 1.0);
   $hold(posedge WCLKN, negedge WADDR[1], 1.0);
   $setup(posedge WADDR[2], posedge WCLKN, 1.0);
   $setup(negedge WADDR[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[2], 1.0);
   $hold(posedge WCLKN, negedge WADDR[2], 1.0);
   $setup(posedge WADDR[3], posedge WCLKN, 1.0);
   $setup(negedge WADDR[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[3], 1.0);
   $hold(posedge WCLKN, negedge WADDR[3], 1.0);
   $setup(posedge WADDR[4], posedge WCLKN, 1.0);
   $setup(negedge WADDR[4], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[4], 1.0);
   $hold(posedge WCLKN, negedge WADDR[4], 1.0);
   $setup(posedge WADDR[5], posedge WCLKN, 1.0);
   $setup(negedge WADDR[5], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[5], 1.0);
   $hold(posedge WCLKN, negedge WADDR[5], 1.0);
   $setup(posedge WADDR[6], posedge WCLKN, 1.0);
   $setup(negedge WADDR[6], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[6], 1.0);
   $hold(posedge WCLKN, negedge WADDR[6], 1.0);
   $setup(posedge WADDR[7], posedge WCLKN, 1.0);
   $setup(negedge WADDR[7], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[7], 1.0);
   $hold(posedge WCLKN, negedge WADDR[7], 1.0);
   $setup(posedge WADDR[8], posedge WCLKN, 1.0);
   $setup(negedge WADDR[8], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[8], 1.0);
   $hold(posedge WCLKN, negedge WADDR[8], 1.0);
   $setup(posedge WADDR[9], posedge WCLKN, 1.0);
   $setup(negedge WADDR[9], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[9], 1.0);
   $hold(posedge WCLKN, negedge WADDR[9], 1.0);
   $setup(posedge WADDR[10], posedge WCLKN, 1.0);
   $setup(negedge WADDR[10], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[10], 1.0);
   $hold(posedge WCLKN, negedge WADDR[10], 1.0);
   $setup(posedge WDATA[0], posedge WCLKN, 1.0);
   $setup(negedge WDATA[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[0], 1.0);
   $hold(posedge WCLKN, negedge WDATA[0], 1.0);
   $setup(posedge WDATA[1], posedge WCLKN, 1.0);
   $setup(negedge WDATA[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[1], 1.0);
   $hold(posedge WCLKN, negedge WDATA[1], 1.0);
   $setup(posedge WCLKE, posedge WCLKN, 1.0);
   $setup(negedge WCLKE, posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WCLKE, 1.0);
   $hold(posedge WCLKN, negedge WCLKE, 1.0);
   $setup(posedge WE, posedge WCLKN, 1.0);
   $setup(negedge WE, posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WE, 1.0);
   $hold(posedge WCLKN, negedge WE, 1.0);
   $setup(posedge RADDR[0], posedge RCLKN, 1.0);
   $setup(negedge RADDR[0], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[0], 1.0);
   $hold(posedge RCLKN, negedge RADDR[0], 1.0);
   $setup(posedge RADDR[1], posedge RCLKN, 1.0);
   $setup(negedge RADDR[1], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[1], 1.0);
   $hold(posedge RCLKN, negedge RADDR[1], 1.0);
   $setup(posedge RADDR[2], posedge RCLKN, 1.0);
   $setup(negedge RADDR[2], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[2], 1.0);
   $hold(posedge RCLKN, negedge RADDR[2], 1.0);
   $setup(posedge RADDR[3], posedge RCLKN, 1.0);
   $setup(negedge RADDR[3], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[3], 1.0);
   $hold(posedge RCLKN, negedge RADDR[3], 1.0);
   $setup(posedge RADDR[4], posedge RCLKN, 1.0);
   $setup(negedge RADDR[4], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[4], 1.0);
   $hold(posedge RCLKN, negedge RADDR[4], 1.0);
   $setup(posedge RADDR[5], posedge RCLKN, 1.0);
   $setup(negedge RADDR[5], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[5], 1.0);
   $hold(posedge RCLKN, negedge RADDR[5], 1.0);
   $setup(posedge RADDR[6], posedge RCLKN, 1.0);
   $setup(negedge RADDR[6], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[6], 1.0);
   $hold(posedge RCLKN, negedge RADDR[6], 1.0);
   $setup(posedge RADDR[7], posedge RCLKN, 1.0);
   $setup(negedge RADDR[7], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[7], 1.0);
   $hold(posedge RCLKN, negedge RADDR[7], 1.0);
   $setup(posedge RADDR[8], posedge RCLKN, 1.0);
   $setup(negedge RADDR[8], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[8], 1.0);
   $hold(posedge RCLKN, negedge RADDR[8], 1.0);
   $setup(posedge RADDR[9], posedge RCLKN, 1.0);
   $setup(negedge RADDR[9], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[9], 1.0);
   $hold(posedge RCLKN, negedge RADDR[9], 1.0);
   $setup(posedge RADDR[10], posedge RCLKN, 1.0);
   $setup(negedge RADDR[10], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[10], 1.0);
   $hold(posedge RCLKN, negedge RADDR[10], 1.0);
   $setup(posedge RCLKE, posedge RCLKN, 1.0);
   $setup(negedge RCLKE, posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RCLKE, 1.0);
   $hold(posedge RCLKN, negedge RCLKE, 1.0);
   $setup(posedge RE, posedge RCLKN, 1.0);
   $setup(negedge RE, posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RE, 1.0);
   $hold(posedge RCLKN, negedge RE, 1.0);
   $recovery(posedge RCLKN, posedge WCLKN, 1.0);
   $recovery(negedge RCLKN, posedge WCLKN, 1.0);
   $removal(posedge RCLKN, posedge WCLKN, 1.0);
   $removal(negedge RCLKN, posedge WCLKN, 1.0);
   $recovery(posedge WCLKN, posedge RCLKN, 1.0);
   $recovery(negedge WCLKN, posedge RCLKN, 1.0);
   $removal(posedge WCLKN, posedge RCLKN, 1.0);
   $removal(negedge WCLKN, posedge RCLKN, 1.0);
endspecify
`endif

endmodule //SB_RAM2048x2NRNW

/*****ice40P08 RAM prims******/

`timescale 10ps/1ps

module SB_IO (
	PACKAGE_PIN, 
	LATCH_INPUT_VALUE, 
	CLOCK_ENABLE, 
	INPUT_CLK, 
	OUTPUT_CLK, 
	OUTPUT_ENABLE, 
	D_OUT_1, 
	D_OUT_0, 
	D_IN_1, 
	D_IN_0
 );

parameter PIN_TYPE			= 6'b000000;	  // The default is set to report IO macros that do not define what IO type is used. 
parameter PULLUP = 1'b0; // by default the IO will have NO pullup, this parameter is used only on bank 0, 1, and 2. Will be ignored when it is placed at bank 3
parameter NEG_TRIGGER = 1'b0; // specify the polarity of all FFs in the IO to be falling edge when NEG_TRIGGER = 1, default is rising edge
parameter IO_STANDARD = "SB_LVCMOS"; // more standards are supported in bank 3 only: SB_SSTL2_CLASS_2, SB_SSTL2_CLASS_1, SB_SSTL18_FULL, SB_SSTL18_HALF
						 // SB_MDDR10, SB_MDDR8, SB_MDDR4, SB_MDDR2

input D_OUT_1;  		// Input output 1
input D_OUT_0;  		// Input output 0

input CLOCK_ENABLE;    		// Clock enables NEW - common to in/out clocks

output D_IN_1;    		// Output input 1
output D_IN_0;    		// Output input 0

input OUTPUT_ENABLE;   		// Ouput-Enable 
input LATCH_INPUT_VALUE;    		// Input control
input INPUT_CLK;   		// Input clock
input OUTPUT_CLK;  		// Output clock

inout 	PACKAGE_PIN; 		//' User's package pin - 'PAD' output

//------------- Main Body of verilog ----------------------------------------------------
wire inclk_, outclk_;
wire inclk, outclk;
reg INCLKE_sync, OUTCLKE_sync; 

assign (weak0, weak1) CLOCK_ENABLE =1'b1 ;
assign inclk_ = (INPUT_CLK ^ NEG_TRIGGER); // change the input clock phase
assign outclk_ = (OUTPUT_CLK ^ NEG_TRIGGER); // change the output clock phase
//assign inclk = (inclk_ & CLOCK_ENABLE);
//assign outclk = (outclk_ & CLOCK_ENABLE);

//////// CLKEN sync ///////
always@(inclk_ or CLOCK_ENABLE)
begin 
    if(~inclk_)
	INCLKE_sync = CLOCK_ENABLE; 
end

always@(outclk_ or CLOCK_ENABLE)
begin 
   if(~outclk_) 	
	OUTCLKE_sync = CLOCK_ENABLE; 
end

assign inclk = (inclk_ & INCLKE_sync);
assign outclk = (outclk_ & OUTCLKE_sync);

wire bs_en;   //Boundary scan enable
wire shift;   //Boundary scan shift
wire tclk;    //Boundary scan clock
wire update;  //Boundary scan update
wire sdi;     //Boundary scan serial data in
wire mode;    //Boundary scan mode
wire hiz_b;   //Boundary scan tristate control
wire sdo;     //Boundary scan serial data out

//wire rstio; disabled as this a power on only signal   	//Normal Input reset
assign  bs_en = 1'b0;	//Boundary scan enable
assign  shift = 1'b0;	//Boundary scan shift
assign  tclk = 1'b0;	//Boundary scan clock
assign  update = 1'b0;	//Boundary scan update
assign  sdi = 1'b0;	//Boundary scan serial data in
assign  mode = 1'b0;	//Boundary scan mode
assign  hiz_b = 1'b1;	//Boundary scan Tristate control
  
wire padoen, padout, padin;
assign PACKAGE_PIN = (~padoen) ? padout : 1'bz;
assign padin = PACKAGE_PIN ;


//parameter Pin_Type  MUST be defined when instantiated
wire hold, oepin;							  // The required package pin type must be set when io_macro is instantiated.
assign hold = LATCH_INPUT_VALUE;
assign oepin = OUTPUT_ENABLE;
 
 preio_physical preiophysical_i (	//original names unchanged
 	.hold(hold),
	.rstio(1'b0),			//Disabled as this is power on only.
	.bs_en(bs_en),
	.shift(shift),
	.tclk(tclk),
	.inclk(inclk),
	.outclk(outclk),
	.update(update),
	.oepin(oepin),
	.sdi(sdi),
	.mode(mode),
	.hiz_b(hiz_b),
	.sdo(sdo),
	.dout1(D_IN_1),
	.dout0(D_IN_0),
	.ddr1(D_OUT_1),
	.ddr0(D_OUT_0),
	.padin(padin),
	.padout(padout),
	.padoen(padoen),
	.cbit(PIN_TYPE)
	);

`ifdef TIMINGCHECK
specify
   (PACKAGE_PIN *> D_IN_0) = (1.0, 1.0);
   (PACKAGE_PIN *> D_IN_1) = (1.0, 1.0);
   (INPUT_CLK *> D_IN_0) = (1.0, 1.0);
   (INPUT_CLK *> D_IN_1) = (1.0, 1.0);
   (D_OUT_0 *> PACKAGE_PIN) = (1.0, 1.0);
   (D_OUT_1 *> PACKAGE_PIN) = (1.0, 1.0);
   (OUTPUT_ENABLE *> PACKAGE_PIN) = (1.0, 1.0);
   (INPUT_CLK *> PACKAGE_PIN) = (1.0, 1.0);
   (OUTPUT_CLK *> PACKAGE_PIN) = (1.0, 1.0);
   (LATCH_INPUT_VALUE *> D_IN_0) = (1.0, 1.0);
   (LATCH_INPUT_VALUE *> D_IN_1) = (1.0, 1.0);
   $setup(posedge CLOCK_ENABLE, posedge INPUT_CLK, 1.0);
   $setup(negedge CLOCK_ENABLE, posedge INPUT_CLK, 1.0);
   $hold(posedge INPUT_CLK, posedge CLOCK_ENABLE, 1.0);
   $hold(posedge INPUT_CLK, negedge CLOCK_ENABLE, 1.0);
   $setup(posedge PACKAGE_PIN, posedge INPUT_CLK, 1.0);
   $setup(negedge PACKAGE_PIN, posedge INPUT_CLK, 1.0);
   $hold(posedge INPUT_CLK, posedge PACKAGE_PIN, 1.0);
   $hold(posedge INPUT_CLK, negedge PACKAGE_PIN, 1.0);
   $setup(posedge PACKAGE_PIN, negedge INPUT_CLK, 1.0);
   $setup(negedge PACKAGE_PIN, negedge INPUT_CLK, 1.0);
   $hold(negedge INPUT_CLK, posedge PACKAGE_PIN, 1.0);
   $hold(negedge INPUT_CLK, negedge PACKAGE_PIN, 1.0);
   $setup(posedge CLOCK_ENABLE, posedge OUTPUT_CLK, 1.0);
   $setup(negedge CLOCK_ENABLE, posedge OUTPUT_CLK, 1.0);
   $hold(posedge OUTPUT_CLK, posedge CLOCK_ENABLE, 1.0);
   $hold(posedge OUTPUT_CLK, negedge CLOCK_ENABLE, 1.0);
   $setup(posedge PACKAGE_PIN, posedge OUTPUT_CLK, 1.0);
   $setup(negedge PACKAGE_PIN, posedge OUTPUT_CLK, 1.0);
   $hold(posedge OUTPUT_CLK, posedge PACKAGE_PIN, 1.0);
   $hold(posedge OUTPUT_CLK, negedge PACKAGE_PIN, 1.0);
   $setup(posedge D_OUT_0, posedge OUTPUT_CLK, 1.0);
   $setup(negedge D_OUT_0, posedge OUTPUT_CLK, 1.0);
   $hold(posedge OUTPUT_CLK, posedge D_OUT_0, 1.0);
   $hold(posedge OUTPUT_CLK, negedge D_OUT_0, 1.0);
   $setup(posedge D_OUT_1, posedge OUTPUT_CLK, 1.0);
   $setup(negedge D_OUT_1, posedge OUTPUT_CLK, 1.0);
   $hold(posedge OUTPUT_CLK, posedge D_OUT_1, 1.0);
   $hold(posedge OUTPUT_CLK, negedge D_OUT_1, 1.0);
   $setup(posedge D_OUT_1, negedge OUTPUT_CLK, 1.0);
   $setup(negedge D_OUT_1, negedge OUTPUT_CLK, 1.0);
   $hold(negedge OUTPUT_CLK, posedge D_OUT_1, 1.0);
   $hold(negedge OUTPUT_CLK, negedge D_OUT_1, 1.0);
   $setup(posedge D_OUT_0, posedge OUTPUT_CLK, 1.0);
   $setup(negedge D_OUT_0, posedge OUTPUT_CLK, 1.0);
   $hold(posedge OUTPUT_CLK, posedge D_OUT_0, 1.0);
   $hold(posedge OUTPUT_CLK, negedge D_OUT_0, 1.0);
   $setup(posedge OUTPUT_ENABLE, posedge OUTPUT_CLK, 1.0);
   $setup(negedge OUTPUT_ENABLE, posedge OUTPUT_CLK, 1.0);
   $hold(posedge OUTPUT_CLK, posedge OUTPUT_ENABLE, 1.0);
   $hold(posedge OUTPUT_CLK, negedge OUTPUT_ENABLE, 1.0);

endspecify
`endif

endmodule

`timescale 10ps/1ps

module SB_GB_IO (
	PACKAGE_PIN, 
	LATCH_INPUT_VALUE, 
	CLOCK_ENABLE, 
	INPUT_CLK, 
	OUTPUT_CLK, 
	OUTPUT_ENABLE, 
	D_OUT_1, 
	D_OUT_0, 
	D_IN_1, 
	D_IN_0,
	GLOBAL_BUFFER_OUTPUT
 );

parameter PIN_TYPE			= 6'b000000;	  // The default is set to report IO macros that do not define what IO type is used. 
parameter PULLUP = 1'b0; // by default the IO will have NO pullup, this parameter is used only on bank 0, 1, and 2. Will be ignored when it is placed at bank 3
parameter NEG_TRIGGER = 1'b0; // specify the polarity of all FFs in the IO to be falling edge when NEG_TRIGGER = 1, default is rising edge
parameter IO_STANDARD = "SB_LVCMOS"; // more standards are supported in bank 3 only: SB_SSTL2_CLASS_2, SB_SSTL2_CLASS_1, SB_SSTL18_FULL, SB_SSTL18_HALF
						 // SB_MDDR10, SB_MDDR8, SB_MDDR4, SB_MDDR2

input D_OUT_1;  		// Input output 1
input D_OUT_0;  		// Input output 0

input CLOCK_ENABLE;    		// Clock enables NEW - common to in/out clocks

output D_IN_1;    		// Output input 1
output D_IN_0;    		// Output input 0

input OUTPUT_ENABLE;   		// Ouput-Enable 
input LATCH_INPUT_VALUE;    		// Input control
input INPUT_CLK;   		// Input clock
input OUTPUT_CLK;  		// Output clock

inout 	PACKAGE_PIN; 		//' User's package pin - 'PAD' output
output GLOBAL_BUFFER_OUTPUT;

//------------- Main Body of verilog ----------------------------------------------------
wire inclk_, outclk_;
wire inclk, outclk;
reg INCLKE_sync,OUTCLKE_sync;

assign (weak0, weak1) CLOCK_ENABLE =1'b1 ;
assign inclk_ = (INPUT_CLK ^ NEG_TRIGGER);
assign outclk_ = (OUTPUT_CLK ^ NEG_TRIGGER);
//assign inclk = (inclk_ & CLOCK_ENABLE);
//assign outclk = (outclk_ & CLOCK_ENABLE);


//////// CLKEN sync ///////
always@(inclk_ or CLOCK_ENABLE)
begin 
    if(~inclk_)
	INCLKE_sync = CLOCK_ENABLE; 
end

always@(outclk_ or CLOCK_ENABLE)
begin 
   if(~outclk_) 	
	OUTCLKE_sync = CLOCK_ENABLE; 
end

assign inclk = (inclk_ & INCLKE_sync);
assign outclk = (outclk_ & OUTCLKE_sync);

wire bs_en;   //Boundary scan enable
wire shift;   //Boundary scan shift
wire tclk;    //Boundary scan clock
wire update;  //Boundary scan update
wire sdi;     //Boundary scan serial data in
wire mode;    //Boundary scan mode
wire hiz_b;   //Boundary scan tristate control
wire sdo;     //Boundary scan serial data out

//wire rstio; disabled as this a power on only signal   	//Normal Input reset

assign  bs_en = 1'b0;	//Boundary scan enable
assign  shift = 1'b0;	//Boundary scan shift
assign  tclk = 1'b0;	//Boundary scan clock
assign  update = 1'b0;	//Boundary scan update
assign  sdi = 1'b0;	//Boundary scan serial data in
assign  mode = 1'b0;	//Boundary scan mode
assign  hiz_b = 1'b1;	//Boundary scan Tristate control
  
wire padoen, padout, padin;
assign PACKAGE_PIN = (~padoen) ? padout : 1'bz;
assign padin = PACKAGE_PIN ;

assign GLOBAL_BUFFER_OUTPUT = padin;


wire hold, oepin;							  // The required package pin type must be set when io_macro is instantiated.
assign hold = LATCH_INPUT_VALUE;
assign oepin = OUTPUT_ENABLE;
 
 preio_physical preiophysical_i (	//original names unchanged
 	.hold(hold),
	.rstio(1'b0),			//Disabled as this is power on only.
	.bs_en(bs_en),
	.shift(shift),
	.tclk(tclk),
	.inclk(inclk),
	.outclk(outclk),
	.update(update),
	.oepin(oepin),
	.sdi(sdi),
	.mode(mode),
	.hiz_b(hiz_b),
	.sdo(sdo),
	.dout1(D_IN_1),
	.dout0(D_IN_0),
	.ddr1(D_OUT_1),
	.ddr0(D_OUT_0),
	.padin(padin),
	.padout(padout),
	.padoen(padoen),
	.cbit(PIN_TYPE)
	);

`ifdef TIMINGCHECK
specify
   (PACKAGE_PIN *> GLOBAL_BUFFER_OUTPUT) = (1.0, 1.0);
   (PACKAGE_PIN *> D_IN_0) = (1.0, 1.0);
   (PACKAGE_PIN *> D_IN_1) = (1.0, 1.0);
   (INPUT_CLK *> D_IN_0) = (1.0, 1.0);
   (INPUT_CLK *> D_IN_1) = (1.0, 1.0);
   (D_OUT_0 *> PACKAGE_PIN) = (1.0, 1.0);
   (D_OUT_1 *> PACKAGE_PIN) = (1.0, 1.0);
   (OUTPUT_ENABLE *> PACKAGE_PIN) = (1.0, 1.0);
   (INPUT_CLK *> PACKAGE_PIN) = (1.0, 1.0);
   (OUTPUT_CLK *> PACKAGE_PIN) = (1.0, 1.0);
   (LATCH_INPUT_VALUE *> D_IN_0) = (1.0, 1.0);
   (LATCH_INPUT_VALUE *> D_IN_1) = (1.0, 1.0);
   $setup(posedge CLOCK_ENABLE, posedge INPUT_CLK, 1.0);
   $setup(negedge CLOCK_ENABLE, posedge INPUT_CLK, 1.0);
   $hold(posedge INPUT_CLK, posedge CLOCK_ENABLE, 1.0);
   $hold(posedge INPUT_CLK, negedge CLOCK_ENABLE, 1.0);
   $setup(posedge PACKAGE_PIN, posedge INPUT_CLK, 1.0);
   $setup(negedge PACKAGE_PIN, posedge INPUT_CLK, 1.0);
   $hold(posedge INPUT_CLK, posedge PACKAGE_PIN, 1.0);
   $hold(posedge INPUT_CLK, negedge PACKAGE_PIN, 1.0);
   $setup(posedge PACKAGE_PIN, negedge INPUT_CLK, 1.0);
   $setup(negedge PACKAGE_PIN, negedge INPUT_CLK, 1.0);
   $hold(negedge INPUT_CLK, posedge PACKAGE_PIN, 1.0);
   $hold(negedge INPUT_CLK, negedge PACKAGE_PIN, 1.0);
   $setup(posedge CLOCK_ENABLE, posedge OUTPUT_CLK, 1.0);
   $setup(negedge CLOCK_ENABLE, posedge OUTPUT_CLK, 1.0);
   $hold(posedge OUTPUT_CLK, posedge CLOCK_ENABLE, 1.0);
   $hold(posedge OUTPUT_CLK, negedge CLOCK_ENABLE, 1.0);
   $setup(posedge PACKAGE_PIN, posedge OUTPUT_CLK, 1.0);
   $setup(negedge PACKAGE_PIN, posedge OUTPUT_CLK, 1.0);
   $hold(posedge OUTPUT_CLK, posedge PACKAGE_PIN, 1.0);
   $hold(posedge OUTPUT_CLK, negedge PACKAGE_PIN, 1.0);
   $setup(posedge D_OUT_0, posedge OUTPUT_CLK, 1.0);
   $setup(negedge D_OUT_0, posedge OUTPUT_CLK, 1.0);
   $hold(posedge OUTPUT_CLK, posedge D_OUT_0, 1.0);
   $hold(posedge OUTPUT_CLK, negedge D_OUT_0, 1.0);
   $setup(posedge D_OUT_1, posedge OUTPUT_CLK, 1.0);
   $setup(negedge D_OUT_1, posedge OUTPUT_CLK, 1.0);
   $hold(posedge OUTPUT_CLK, posedge D_OUT_1, 1.0);
   $hold(posedge OUTPUT_CLK, negedge D_OUT_1, 1.0);
   $setup(posedge D_OUT_1, negedge OUTPUT_CLK, 1.0);
   $setup(negedge D_OUT_1, negedge OUTPUT_CLK, 1.0);
   $hold(negedge OUTPUT_CLK, posedge D_OUT_1, 1.0);
   $hold(negedge OUTPUT_CLK, negedge D_OUT_1, 1.0);
   $setup(posedge D_OUT_0, posedge OUTPUT_CLK, 1.0);
   $setup(negedge D_OUT_0, posedge OUTPUT_CLK, 1.0);
   $hold(posedge OUTPUT_CLK, posedge D_OUT_0, 1.0);
   $hold(posedge OUTPUT_CLK, negedge D_OUT_0, 1.0);
   $setup(posedge OUTPUT_ENABLE, posedge OUTPUT_CLK, 1.0);
   $setup(negedge OUTPUT_ENABLE, posedge OUTPUT_CLK, 1.0);
   $hold(posedge OUTPUT_CLK, posedge OUTPUT_ENABLE, 1.0);
   $hold(posedge OUTPUT_CLK, negedge OUTPUT_ENABLE, 1.0);

endspecify
`endif

endmodule



`timescale 1ps/1ps
module SB_GB (	
GLOBAL_BUFFER_OUTPUT,
USER_SIGNAL_TO_GLOBAL_BUFFER);

input USER_SIGNAL_TO_GLOBAL_BUFFER;			
output GLOBAL_BUFFER_OUTPUT;	

assign GLOBAL_BUFFER_OUTPUT = USER_SIGNAL_TO_GLOBAL_BUFFER;

`ifdef TIMINGCHECK
specify
   (USER_SIGNAL_TO_GLOBAL_BUFFER *> GLOBAL_BUFFER_OUTPUT) = (1.0, 1.0);
endspecify
`endif


endmodule	//SB_GB


`timescale 10ps/1ps


//************************************************

//************************************************


`timescale 1ps/1ps
module preio_physical 	(hold, rstio, bs_en, shift, tclk, inclk, outclk, update, oepin, sdi, mode, 
			hiz_b, sdo, dout1, dout0, ddr1, ddr0, padin, padout, padoen, cbit);

input bs_en;   //JTAG enable
input shift;   //JTAG shift
input tclk;    //JTAG clock
input update;  //JTAG update
input sdi;     //JTAG serial data in
input mode;    //JTAG mode
input hiz_b;   //JTAG high X control
output sdo;    //JTAG serial data out

output dout1;  //Normal Input cell output 1
output dout0;  //Normal Input cell output 0
input ddr1;    //Normal Output cell input 1
input ddr0;    //Normal Output cell input 0
input oepin;   //Normal Ouput-Enable 
input hold;    //Normal Input cell control
input rstio;   //Normal Input cell reset
input inclk;   //Normal Input cell clock
input outclk;  //Normal Output cell clock

input [5:0] cbit; //Configurion bits

input 	padin;   //PAD input
output 	padout;  //PAD output
output	padoen;  //PAD output enable




//Signals declaration
wire padin_n1;
wire inclk_n2;
wire padin_n3;
reg  in_MUX_n4 = 0;
wire hold_AND2;
wire dout0;

wire ddr0_n11;
wire outclk_n12;
wire ddr1_n13;
wire n14;
wire dout_reg_0_n;

wire Reg_or_Wire_N17;
wire n18;
//wire n19;
reg n19; 

wire tristate;
wire outclk_n22;
wire n26;

reg  oen_n_n24 = 0;
wire jtag_update_n30;

reg din_reg_0 = 0;
reg din_reg_1 = 0;
reg dout_reg_0 = 0;
reg dout_reg_1 = 0;
reg tristate_q = 0;
reg jtag_oe_reg = 0;

					
// Miscc logics
//---------------------

assign jtag_update_n30 = ~( bs_en & (~update ) );

//---------------------------------------------------------------------------
//
//	Assign output
//
//---------------------------------------------------------------------------
assign sdo = din_reg_0;
assign dout1 = din_reg_1;

//---------------------------------------------------------------------------
//
//	Input logic
//
//---------------------------------------------------------------------------

assign padin_n1 = (shift) ? dout_reg_0  : padin;

assign inclk_n2 = (bs_en) ? tclk : inclk;

always @(posedge inclk_n2 or posedge rstio)
   if (rstio) din_reg_0 <= 1'b0 ; //#1 1'b0;
   else din_reg_0 <= padin_n1;    //#1 padin_n1;

assign padin_n3 = (bs_en) ? din_reg_0 : padin;

always @(negedge inclk_n2 or posedge rstio)
   if (rstio) din_reg_1 <= 1'b0 ; // #1 1'b0;
   else if (jtag_update_n30) din_reg_1 <= padin_n3; //  #1 padin_n3;

assign hold_AND2 = cbit[1] & hold;

// 	Input MUX
always @(hold_AND2, cbit[0], dout0, padin, din_reg_0) begin 
   case ({hold_AND2, cbit[0]})
      2'b00 : 	in_MUX_n4 = din_reg_0;
      2'b01 : 	in_MUX_n4 = padin;
      2'b10 : 	in_MUX_n4 = dout0;
      2'b11 : 	in_MUX_n4 = dout0;
      default : in_MUX_n4 = 1'b0;
      endcase
 end     
 
assign dout0 = (mode) ? din_reg_1 : in_MUX_n4;


// Output Register
always @(posedge outclk_n12 or posedge rstio)
   if (rstio) dout_reg_0 <=  1'b0 ; //#1 1'b0;
   else dout_reg_0 <=  ddr0_n11 ; // #1 ddr0_n11;

// Muxes for Output registers
assign dout_reg_0_n = ~dout_reg_0;
assign Reg_or_Wire_N17 = cbit[2] ? dout_reg_0_n : ddr0;
assign n18 = n19 ? dout_reg_1 : dout_reg_0;
//assign n19 = ~(outclk_n12 || cbit[2]);

always@(outclk_n12,cbit[2])
begin 
	n19<= ~(outclk_n12 || cbit[2]);
end 


assign n14 = cbit[3] ? Reg_or_Wire_N17 : n18;
assign padout = mode ? dout_reg_1 : n14;

// JTAG Assigns
assign ddr0_n11 = (shift) ? tristate_q  : ddr0;

assign outclk_n12 = (bs_en) ? tclk : outclk;
assign ddr1_n13 = (bs_en) ? dout_reg_0 : ddr1;

// JTAG register 
always @(negedge outclk_n12 or posedge rstio)
   if (rstio) dout_reg_1 <=  1'b0 ; //#1 1'b0;
   else if (jtag_update_n30) dout_reg_1 <= ddr1_n13; //  #1 ddr1_n13;

//---------------------------------------------------------------------------
//
//	Output Enable Logic
//
//---------------------------------------------------------------------------

// OE Tristate Register
assign tristate = (shift) ? sdi  : oepin;
always @(posedge outclk_n22 or posedge rstio)
   if (rstio) tristate_q <= 1'b0;	// #1 1'b0;
   else tristate_q <= tristate;

// JTAG register
assign outclk_n22 = (bs_en) ? tclk : outclk;
always @(negedge outclk_n22 or posedge rstio)
   if (rstio) jtag_oe_reg <=  1'b0 ; // #1 1'b0;
   else if (jtag_update_n30) jtag_oe_reg <= padin_n3;

always @(cbit[5],cbit[4], oepin, tristate_q)  begin 
   case ({cbit[5],cbit[4]})
      2'b00 : oen_n_n24 = 1'b0;
      2'b01 : oen_n_n24 = 1'b1;
      2'b10 : oen_n_n24 = oepin;
      2'b11 : oen_n_n24 = tristate_q;
 
   endcase
end      
		

assign n26 = (mode) ? jtag_oe_reg : oen_n_n24;

assign padoen = ~(hiz_b & n26);

endmodule //preio_physical


// Warm boot, {s1, s0} used to select one of the four boot addresses
// s1 s0  boot_addr
// 0  0   0
// 0  1   1
// 1  0   2
// 1  1   3

`timescale 1ps/1ps
module SB_WARMBOOT (	
BOOT, S1, S0);

input BOOT, S1, S0;			

endmodule	//SB_WARMBOOT

`timescale 1ps/1ps
// Differential signaling IO
module SB_IO_DS (
	PACKAGE_PIN, 
	PACKAGE_PIN_B, 
	LATCH_INPUT_VALUE, 
	CLOCK_ENABLE, 
	INPUT_CLK, 
	OUTPUT_CLK, 
	OUTPUT_ENABLE, 
	D_OUT_1, 
	D_OUT_0, 
	D_IN_1, 
	D_IN_0
 );

parameter PIN_TYPE			= 6'b000000;	  // The default is set to report IO macros that do not define what IO type is used. 
parameter NEG_TRIGGER = 1'b0; // specify the polarity of all FFs in the IO to be falling edge when NEG_TRIGGER = 1, default is rising edge
parameter IO_STANDARD = "SB_LVDS_OUTPUT"; // another supported standard is SB_LVDS_IO 

input D_OUT_1;  		// Input output 1
input D_OUT_0;  		// Input output 0

input CLOCK_ENABLE;    		// Clock enables NEW - common to in/out clocks

output D_IN_1;    		// Output input 1
output D_IN_0;    		// Output input 0

input OUTPUT_ENABLE;   		// Ouput-Enable 
input LATCH_INPUT_VALUE;    		// Input control
input INPUT_CLK;   		// Input clock
input OUTPUT_CLK;  		// Output clock

inout 	PACKAGE_PIN; 		//' User's package pin - 'PAD' output
inout 	PACKAGE_PIN_B; 		//' User's package pin - 'PAD' output


//------------- Main Body of verilog ----------------------------------------------------
wire inclk_, outclk_;
wire inclk, outclk;
reg INCLKE_sync,OUTCLKE_sync;

assign (weak0, weak1) CLOCK_ENABLE =1'b1 ;
assign inclk_ = (INPUT_CLK ^ NEG_TRIGGER); // change the input clock phase
assign outclk_ = (OUTPUT_CLK ^ NEG_TRIGGER); // change the output clock phase
//assign inclk = (inclk_ & CLOCK_ENABLE);
//assign outclk = (outclk_ & CLOCK_ENABLE);


//////// CLKEN sync ///////
always@(inclk_ or CLOCK_ENABLE)
begin 
    if(~inclk_)
	INCLKE_sync = CLOCK_ENABLE; 
end

always@(outclk_ or CLOCK_ENABLE)
begin 
   if(~outclk_) 	
	OUTCLKE_sync = CLOCK_ENABLE; 
end

assign inclk = (inclk_ & INCLKE_sync);
assign outclk = (outclk_ & OUTCLKE_sync);

wire bs_en;   //Boundary scan enable
wire shift;   //Boundary scan shift
wire tclk;    //Boundary scan clock
wire update;  //Boundary scan update
wire sdi;     //Boundary scan serial data in
wire mode;    //Boundary scan mode
wire hiz_b;   //Boundary scan tristate control
wire sdo;     //Boundary scan serial data out

//wire rstio; disabled as this a power on only signal   	//Normal Input reset

assign  bs_en = 1'b0;	//Boundary scan enable
assign  shift = 1'b0;	//Boundary scan shift
assign  tclk = 1'b0;	//Boundary scan clock
assign  update = 1'b0;	//Boundary scan update
assign  sdi = 1'b0;	//Boundary scan serial data in
assign  mode = 1'b0;	//Boundary scan mode
assign  hiz_b = 1'b1;	//Boundary scan Tristate control
  
wire padoen, padout, padin;
assign PACKAGE_PIN = (~padoen) ? padout : 1'bz;
assign PACKAGE_PIN_B = (~padoen) ? ~padout : 1'bz;

assign padin = PACKAGE_PIN ;


//parameter Pin_Type  MUST be defined when instantiated
wire hold, oepin;							  // The required package pin type must be set when io_macro is instantiated.
assign hold = LATCH_INPUT_VALUE;
assign oepin = OUTPUT_ENABLE;
 
 preio_physical preiophysical_i (	//original names unchanged
 	.hold(hold),
	.rstio(1'b0),			//Disabled as this is power on only.
	.bs_en(bs_en),
	.shift(shift),
	.tclk(tclk),
	.inclk(inclk),
	.outclk(outclk),
	.update(update),
	.oepin(oepin),
	.sdi(sdi),
	.mode(mode),
	.hiz_b(hiz_b),
	.sdo(sdo),
	.dout1(D_IN_1),
	.dout0(D_IN_0),
	.ddr1(D_OUT_1),
	.ddr0(D_OUT_0),
	.padin(padin),
	.padout(padout),
	.padoen(padoen),
	.cbit(PIN_TYPE)
	);

`ifdef TIMINGCHECK
specify
   (PACKAGE_PIN *> D_IN_0) = (1.0, 1.0);
   (PACKAGE_PIN_B *> D_IN_0) = (1.0, 1.0);
   (INPUT_CLK *> D_IN_0) = (1.0, 1.0);
   (INPUT_CLK *> D_IN_1) = (1.0, 1.0);
   (INPUT_CLK *> PACKAGE_PIN) = (1.0, 1.0);
   (INPUT_CLK *> PACKAGE_PIN_B) = (1.0, 1.0);
   (D_OUT_0 *> PACKAGE_PIN) = (1.0, 1.0);
   (D_OUT_0 *> PACKAGE_PIN_B) = (1.0, 1.0);
   (D_OUT_1 *> PACKAGE_PIN) = (1.0, 1.0);
   (D_OUT_1 *> PACKAGE_PIN_B) = (1.0, 1.0);
   (OUTPUT_ENABLE *> PACKAGE_PIN) = (1.0, 1.0);
   (OUTPUT_ENABLE *> PACKAGE_PIN_B) = (1.0, 1.0);
   (LATCH_INPUT_VALUE *> D_IN_0) = (1.0, 1.0);
   (LATCH_INPUT_VALUE *> D_IN_1) = (1.0, 1.0);
   (OUTPUT_CLK *> PACKAGE_PIN) = (1.0, 1.0);
   (OUTPUT_CLK *> PACKAGE_PIN_B) = (1.0, 1.0);

   $setup(posedge CLOCK_ENABLE, posedge INPUT_CLK, 1.0);
   $setup(negedge CLOCK_ENABLE, posedge INPUT_CLK, 1.0);
   $hold(posedge INPUT_CLK, posedge CLOCK_ENABLE, 1.0);
   $hold(posedge INPUT_CLK, negedge CLOCK_ENABLE, 1.0);
   $setup(posedge PACKAGE_PIN, posedge INPUT_CLK, 1.0);
   $setup(negedge PACKAGE_PIN, posedge INPUT_CLK, 1.0);
   $setup(posedge PACKAGE_PIN_B, posedge INPUT_CLK, 1.0);
   $setup(negedge PACKAGE_PIN_B, posedge INPUT_CLK, 1.0);
   $hold(posedge INPUT_CLK, posedge PACKAGE_PIN, 1.0);
   $hold(posedge INPUT_CLK, negedge PACKAGE_PIN, 1.0);
   $hold(posedge INPUT_CLK, posedge PACKAGE_PIN_B, 1.0);
   $hold(posedge INPUT_CLK, negedge PACKAGE_PIN_B, 1.0);
   $setup(posedge PACKAGE_PIN, negedge INPUT_CLK, 1.0);
   $setup(negedge PACKAGE_PIN, negedge INPUT_CLK, 1.0);
   $hold(negedge INPUT_CLK, posedge PACKAGE_PIN, 1.0);
   $hold(negedge INPUT_CLK, negedge PACKAGE_PIN, 1.0);
   $setup(posedge PACKAGE_PIN_B, negedge INPUT_CLK, 1.0);
   $setup(negedge PACKAGE_PIN_B, negedge INPUT_CLK, 1.0);
   $hold(negedge INPUT_CLK, posedge PACKAGE_PIN_B, 1.0);
   $hold(negedge INPUT_CLK, negedge PACKAGE_PIN_B, 1.0);
   $setup(posedge CLOCK_ENABLE, posedge OUTPUT_CLK, 1.0);
   $setup(negedge CLOCK_ENABLE, posedge OUTPUT_CLK, 1.0);
   $hold(posedge OUTPUT_CLK, posedge CLOCK_ENABLE, 1.0);
   $hold(posedge OUTPUT_CLK, negedge CLOCK_ENABLE, 1.0);
   $setup(posedge PACKAGE_PIN, posedge OUTPUT_CLK, 1.0);
   $setup(negedge PACKAGE_PIN, posedge OUTPUT_CLK, 1.0);
   $hold(posedge OUTPUT_CLK, posedge PACKAGE_PIN, 1.0);
   $hold(posedge OUTPUT_CLK, negedge PACKAGE_PIN, 1.0);
   $setup(posedge PACKAGE_PIN_B, posedge OUTPUT_CLK, 1.0);
   $setup(negedge PACKAGE_PIN_B, posedge OUTPUT_CLK, 1.0);
   $hold(posedge OUTPUT_CLK, posedge PACKAGE_PIN_B, 1.0);
   $hold(posedge OUTPUT_CLK, negedge PACKAGE_PIN_B, 1.0);
   $setup(posedge D_OUT_0, posedge OUTPUT_CLK, 1.0);
   $setup(negedge D_OUT_0, posedge OUTPUT_CLK, 1.0);
   $hold(posedge OUTPUT_CLK, posedge D_OUT_0, 1.0);
   $hold(posedge OUTPUT_CLK, negedge D_OUT_0, 1.0);
   $setup(posedge D_OUT_1, posedge OUTPUT_CLK, 1.0);
   $setup(negedge D_OUT_1, posedge OUTPUT_CLK, 1.0);
   $hold(posedge OUTPUT_CLK, posedge D_OUT_1, 1.0);
   $hold(posedge OUTPUT_CLK, negedge D_OUT_1, 1.0);
   $setup(posedge D_OUT_1, negedge OUTPUT_CLK, 1.0);
   $setup(negedge D_OUT_1, negedge OUTPUT_CLK, 1.0);
   $hold(negedge OUTPUT_CLK, posedge D_OUT_1, 1.0);
   $hold(negedge OUTPUT_CLK, negedge D_OUT_1, 1.0);
   $setup(posedge D_OUT_0, posedge OUTPUT_CLK, 1.0);
   $setup(negedge D_OUT_0, posedge OUTPUT_CLK, 1.0);
   $hold(posedge OUTPUT_CLK, posedge D_OUT_0, 1.0);
   $hold(posedge OUTPUT_CLK, negedge D_OUT_0, 1.0);
   $setup(posedge OUTPUT_ENABLE, posedge OUTPUT_CLK, 1.0);
   $setup(negedge OUTPUT_ENABLE, posedge OUTPUT_CLK, 1.0);
   $hold(posedge OUTPUT_CLK, posedge OUTPUT_ENABLE, 1.0);
   $hold(posedge OUTPUT_CLK, negedge OUTPUT_ENABLE, 1.0);

endspecify
`endif

endmodule


`timescale 1ps/1ps
module GND (Y);

    output Y;
supply0 Y ;
endmodule


`timescale 1ps/1ps
module VCC(Y);

    output Y;

supply1 Y ;

endmodule

/****PLL Primitives****/

`timescale 1ps/1ps

module ShiftReg (clk, init, phase0, phase90, phase180, phase270);
input clk, init; 
output phase0, phase90, phase180, phase270;

reg phase0, phase90, phase180, phase270;

always @ (posedge clk or posedge init)
   begin
	if (init)  
		begin
			phase0	 = 1'b0;
			phase90  = 1'b0;
			phase180 = 1'b1;
			phase270 = 1'b1;
		end
	else	
		begin
   	    	phase0 	 <=	phase270;
   	    	phase90  <=	phase0;
   	    	phase180 <=	phase90;
   	    	phase270 <=	phase180;
		end
    end
endmodule

/*
module mux2to1 (a, b, select, out); 
  input a,b; 
  input select; 
  output out; 
  reg    out;
 
  always @ (a or b or select) 
  begin 
    case (select) 
      1'b0   : out = a; 
      1'b1   : out = b; 
    endcase 
  end 

endmodule //mux2to1
*/

/*
`timescale 1ps/1ps
module mux4to1 (a, b, c, d, select, o); 
  input a,b,c,d; 
  input  [1:0] select; 
  output o; 
  reg    o;
 
  always @ (a or b or c or d or select) 
  begin 
    case (select) 
      2'b00   : o = a; 
      2'b01   : o = b; 
      2'b10   : o = c; 
      2'b11	  : o = d; 
    endcase 
  end 

endmodule //mux4to1
*/ 

/*
`timescale 1ps/1ps
module FineDlyAdj ( DlyAdj, signalin, delayedout);
	input signalin;
	input [3:0] DlyAdj;
	output delayedout;
	parameter FIXED_DELAY_ADJUSTMENT = 4'b0000;
	parameter DELAY_ADJUSTMENT_MODE = "FIXED";
	reg test_signalin;
	reg delayedout;

	integer buf_delay = 150;  //In picoseconds
	integer non_variable_delay = 100;
	integer num_bufs = 0;
	integer total_delay;
	wire [3:0] fixed_delay_adj = FIXED_DELAY_ADJUSTMENT;
	
	wire [3:0] bufcntselector = (DELAY_ADJUSTMENT_MODE == "DYNAMIC") ? DlyAdj : fixed_delay_adj;

initial
begin
    if (DELAY_ADJUSTMENT_MODE == "FIXED" && (FIXED_DELAY_ADJUSTMENT > 15 || FIXED_DELAY_ADJUSTMENT < 0))
       begin
	     $display ("************************SBT: Error****************************");
	     $display ("Valid values for FIXED_DELAY_ADJUSTMENT parameter are 0 - 15");
	     $display ("**************************************************************");
	     $finish;
	    end
	  if ((DELAY_ADJUSTMENT_MODE == "DYNAMIC" && FIXED_DELAY_ADJUSTMENT != 0))
	    begin
	     $display ("************************SBT: Info*****************************");
	     $display ("Since DELAY_ADJUSTMENT_MODE=\"DYNAMIC\", parameter FIXED_DELAY_ADJUSTMENT will be ignored.");
		 $display ("Set FIXED_DELAY_ADJUSTMENT=0 to disable this message.");
	     $display ("**************************************************************");
	    end
end

 always @ (signalin or bufcntselector) 
  begin 
    case (bufcntselector) 
      4'b0000   : num_bufs = 1; 
      4'b0001   : num_bufs = 2; 
      4'b0010   : num_bufs = 3; 
      4'b0011   : num_bufs = 4; 
      4'b0100   : num_bufs = 5; 
      4'b0101   : num_bufs = 6; 
      4'b0110   : num_bufs = 7; 
      4'b0111   : num_bufs = 8; 
      4'b1000   : num_bufs = 9; 
      4'b1001   : num_bufs = 10; 
      4'b1010   : num_bufs = 11; 
      4'b1011   : num_bufs = 12; 
      4'b1100   : num_bufs = 13; 
      4'b1101   : num_bufs = 14; 
      4'b1110   : num_bufs = 15; 
      4'b1111   : num_bufs = 16; 
      default   :  begin       
	     $display ("************************SBT: Attention************************");
	     $display ("Fine Delay Adjustment Values have not been specified correctly.");
	     $display ("If you wish to control the delay dynamically, please check that the DYNAMICDELAY port is connected and DELAY_ADJUSTMENT_MODE = \"DYNAMIC\"");
	     $display ("If you wish to wish to set a fixed delay, please specify DELAY_ADJUSTMENT_MODE = \"FIXED\" and the delay value using the FIXED_DELAY_ADJUSTMENT parameter.");
	     $display ("**************************************************************");
	            end

    endcase 
  
   total_delay = non_variable_delay + (num_bufs*buf_delay);
   # total_delay;
   delayedout <= signalin;
  
end 
 
endmodule	//FineDlyAdj
*/
/* 

`timescale 1ps/1ps
module Delay4Buf (a, s, delay4bufout, muxinvout);
input a;
input [1:0] s;
output delay4bufout, muxinvout;
parameter BUF_DELAY = 150;
parameter MUXINV_DELAY = 100; 

buf # BUF_DELAY  bufinst1 (buf1out, a);
buf # BUF_DELAY  bufinst2 (buf2out, buf1out);
buf # BUF_DELAY  bufinst3 (buf3out, buf2out);
buf # BUF_DELAY  bufinst4 (delay4bufout, buf3out);


mux4to1 muxinst (.a(buf1out), .b(buf2out), .c(buf3out), .d(delay4bufout), .select(s), .o(muxout));
not # MUXINV_DELAY (muxinvout, muxout);

endmodule
*/ 

/*

`timescale 1ps/1ps
module FineDlyAdj (DlyAdj, signalin, delayedout);
	input signalin;
	input [3:0] DlyAdj;
	output delayedout;
	parameter FIXED_DELAY_ADJUSTMENT = 4'b0000;
	parameter DELAY_ADJUSTMENT_MODE = "FIXED";
	wire delayedout;
	wire l2muxout;

	parameter BUF_DELAY = 150;
	parameter MUXINV_DELAY = 0; //100; Modified to make consistent with STA

wire [3:0] fixed_delay_adj = FIXED_DELAY_ADJUSTMENT;
wire [3:0] bufcntselector = (DELAY_ADJUSTMENT_MODE == "DYNAMIC")? DlyAdj : fixed_delay_adj;

initial
begin
  if (DELAY_ADJUSTMENT_MODE == "FIXED" && (FIXED_DELAY_ADJUSTMENT > 15 || FIXED_DELAY_ADJUSTMENT < 0))
     begin
	    $display ("************************SBT: ERROR ****************************");
	    $display ("Valid values for FIXED_DELAY_ADJUSTMENT parameter are 4'b0000 through 4'b1111");
	    $display ("Due to incorrect configuration of the PLL, the simulation results are invalid.");
	    $display ("**************************************************************");
	    $display ("Exiting simulation");
	    $finish;
	 end
    if ((DELAY_ADJUSTMENT_MODE == "DYNAMIC" && FIXED_DELAY_ADJUSTMENT != 0))
	 begin
	    $display ("************************SBT: Info*****************************");
	    $display ("Since DELAY_ADJUSTMENT_MODE=\"DYNAMIC\", parameter FIXED_DELAY_ADJUSTMENT will be ignored.");
	    $display ("Set FIXED_DELAY_ADJUSTMENT=0 to disable this message.");
	    $display ("**************************************************************");
	 end
end

Delay4Buf delay4bufinst1 (.a(signalin), .s(bufcntselector[1:0]), .delay4bufout(delay4bufout1), .muxinvout(muxinvout1));
defparam delay4bufinst1.BUF_DELAY = BUF_DELAY;
defparam delay4bufinst1.MUXINV_DELAY = MUXINV_DELAY;

Delay4Buf delay4bufinst2 (.a(delay4bufout1), .s(bufcntselector[1:0]), .delay4bufout(delay4bufout2), .muxinvout(muxinvout2));
defparam delay4bufinst2.BUF_DELAY = BUF_DELAY;
defparam delay4bufinst2.MUXINV_DELAY = MUXINV_DELAY;

Delay4Buf delay4bufinst3 (.a(delay4bufout2), .s(bufcntselector[1:0]), .delay4bufout(delay4bufout3), .muxinvout(muxinvout3));
defparam delay4bufinst3.BUF_DELAY = BUF_DELAY;
defparam delay4bufinst3.MUXINV_DELAY = MUXINV_DELAY;

Delay4Buf delay4bufinst4 (.a(delay4bufout3), .s(bufcntselector[1:0]), .delay4bufout(delay4bufout4), .muxinvout(muxinvout4));
defparam delay4bufinst4.BUF_DELAY = BUF_DELAY;
defparam delay4bufinst4.MUXINV_DELAY = MUXINV_DELAY;

mux4to1 level2muxinst (.a(muxinvout1), .b(muxinvout2), .c(muxinvout3), .d(muxinvout4), .select(bufcntselector[3:2]), .o(l2muxout));
not # MUXINV_DELAY level2invinst(delayedout, l2muxout);

endmodule	//FineDlyAdj
*/ 



`timescale 1ps/1ps	
module SbtSPLL (
		REFERENCECLK,
		EXTFEEDBACK,
		DYNAMICDELAY,
		BYPASS,	
		RESET,		
		
		PLLOUT,		
		LOCK   		
);

//----------------------------------------------------------------------
// Port Declarations
//----------------------------------------------------------------------

// Inputs

input REFERENCECLK;		//Driven by core logic
input	EXTFEEDBACK;  			//Driven by core logic
input	[3:0] DYNAMICDELAY;  	//Driven by core logic
input	BYPASS;				//Driven by core logic
input	RESET;				//Driven by core logic

// Outputs
output 	PLLOUT;		//PLL output to core logic
output	LOCK;				//Output of PLL

//Frequency Specification
//parameter REFERENCE_CLK_FREQUENCY = 100; 		//Floating Point
//parameter PLLOUT_FREQUENCY = 100;			//Floating Point

//Feedback
parameter FEEDBACK_PATH = "SIMPLE";	//String  (simple, delay, phase_and_delay, external) (3 cbits, not 2)
			// If "external" check for signal connectivity on EXTFEEDBACK port.
parameter DELAY_ADJUSTMENT_MODE = "NONE"; //String. If FEEDBACK_SELECT="external",
				// specify DELAY_ADJUSTMENT_MODE as DYNAMIC or FIXED 
				// Check for signal connectivity on DYNAMIC_DELAY[3:0] 
				// && EXTFEEDBACK port
parameter FIXED_DELAY_ADJUSTMENT = 4'b0000; 		//Integer. Specify only if 
				//FEEDBACK_SELECT_MODE="external" && DELAY_ADJUSTMENT_MODE = "fixed". 

//Phase shifted or direct output (3 cbits)
parameter PLLOUT_PHASE = "NONE"; //0deg,90deg,180deg,270deg,none

//Use the Spreadsheet to populate the values below.
parameter DIVR = 4'b0000; 	//determine a good default value
parameter DIVF = 6'b000000; //determine a good default value
parameter DIVQ = 3'b000; 	//determine a good default value
parameter FILTER_RANGE = 3'b000; 	//determine a good default value

//Additional cbits
parameter ENABLE_ICEGATE = 1'b0;

wire ABPLLOUT;
wire phaseShiftMuxOutNet;
wire FSEnet;
wire FBnet;
wire finedelayin, finedelayout;
wire [5:0] DIVFBus = DIVF; 
wire [3:0] DIVRBus = DIVR; 
wire [2:0] DIVQBus = DIVQ; 
wire [2:0] RANGEBus = FILTER_RANGE; 

reg [1:0] phasesel;
reg [1:0] delaymuxsel;
//reg fbout;

initial
begin
 if (PLLOUT_PHASE == "0deg")
    phasesel = 2'b00;
else if (PLLOUT_PHASE == "90deg")
    phasesel = 2'b01;
else if (PLLOUT_PHASE == "180deg")
    phasesel = 2'b10;
else if (PLLOUT_PHASE == "270deg")
    phasesel = 2'b11;
else if (PLLOUT_PHASE != "NONE")
   begin
	        $display ("************************SBT : ERROR ****************************");
	        $display ("Parameter PLLOUT_PHASE is set to an illegal value.");
	        $display ("Legal values should be one of \"NONE\", \"0deg\", \"90deg\", \"180deg\", \"270deg\". ");
	        $display ("Due to incorrect configuration of the PLL, the simulation results are invalid.");
	        $display ("***************************************************************");
	        $finish;
   end
end


assign PLLOUT = (BYPASS == 1'b1) ? REFERENCECLK : ((PLLOUT_PHASE == "NONE") ? ABPLLOUT : phaseShiftMuxOutNet);
assign FSEnet = (FEEDBACK_PATH == "SIMPLE") ? 1'b1 : 1'b0;
assign FBnet = (FEEDBACK_PATH == "SIMPLE") ? 1'b0 : finedelayout;


initial
begin

 if (FEEDBACK_PATH != "EXTERNAL")
 	begin
	    $display ("************************SBT : Info*****************************");
	    $display ("Note that any signal connection to the EXTFEEDBACK port of the PLL will be ignored");
	    $display ("***************************************************************");
	   	end
 if (FEEDBACK_PATH == "EXTERNAL")
    begin 
       delaymuxsel = 2'b11;
        if ( (DELAY_ADJUSTMENT_MODE != "FIXED") && (DELAY_ADJUSTMENT_MODE != "DYNAMIC") )
		begin
	        $display ("************************SBT : ERROR ************************");
	        $display ("Since FEEDBACK_PATH=\"EXTERNAL\", DELAY_ADJUSTMENT_MODE should be \"FIXED\" or \"DYNAMIC\"");
	        $display ("Due to incorrect configuration of the PLL, the simulation results are invalid.");
	        $display ("***************************************************************");
	        $finish;
		end
		if (PLLOUT_PHASE != "NONE")
		begin
	        $display ("************************ SBT : ERROR **************************");
	        $display ("Since FEEDBACK_PATH=\"EXTERNAL\", Phase Adjustment is NOT permitted. Please set PLLOUT_PHASE=\"NONE\"");
	        $display ("*************************************************************");
	        $finish;
		end
    end				
 else if (FEEDBACK_PATH == "DELAY")
    begin 
    	delaymuxsel = 2'b00;
        if ( (DELAY_ADJUSTMENT_MODE != "FIXED") && (DELAY_ADJUSTMENT_MODE != "DYNAMIC") )
		begin
	        $display ("************************ SBT : ERROR **************************");
	        $display ("Since FEEDBACK_PATH=\"DELAY\", DELAY_ADJUSTMENT_MODE should be \"FIXED\" or \"DYNAMIC\"");
	        $display ("Due to incorrect configuration of the PLL, the simulation results are invalid.");
	        $display ("***************************************************************");
	        $finish;
		end
		if (PLLOUT_PHASE != "NONE")
		begin 
	        $display ("************************ SBT : ERROR **************************");
	        $display ("Since FEEDBACK_PATH=\"DELAY\", Phase Adjustment is NOT permitted. Please set PLLOUT_PHASE=\"NONE\"");
		     $display ("Due to incorrect configuration of the PLL, the simulation results are invalid.");
	        $display ("***************************************************************");
	        $finish;
		end
    end				
 else if (FEEDBACK_PATH == "PHASE_AND_DELAY")
	begin
    	delaymuxsel = 2'b01;
        if ( (DELAY_ADJUSTMENT_MODE != "FIXED") && (DELAY_ADJUSTMENT_MODE != "DYNAMIC") )
		begin
	        $display ("************************SBT : Attention************************");
	        $display ("Since FEEDBACK_PATH=\"PHASE_AND_DELAY\", DELAY_ADJUSTMENT_MODE should be FIXED or DYNAMIC");
	        $display ("***************************************************************");
		end
		if ( (PLLOUT_PHASE != "0deg") && (PLLOUT_PHASE != "90deg" )
				&& (PLLOUT_PHASE != "180deg") && (PLLOUT_PHASE != "270deg") )
		begin
	        $display ("************************SBT : Attention************************");
	        $display ("FEEDBACK_PATH=\"PHASE_AND_DELAY\", but PLLOUT_PHASE is not specified correctly");
	        $display ("***************************************************************");
		end
    end				
else if (FEEDBACK_PATH == "SIMPLE")
   begin
		//Ignore DELAY_ADJUSTMENT_MODE, FIXED_DELAY_ADJUSTMENT   
	  $display ("************************SBT : Attention***************************");
	  $display ("Since FEEDBACK_PATH=\"SIMPLE\", the FIXED_DELAY_ADJUSTMENT value will be ignored");
	  $display ("******************************************************************");


    if (PLLOUT_PHASE != "NONE")
		begin
	        $display ("************************SBT : Attention***************************");
	        $display ("The PLL output frequency will be divided by 4 and phase shifted.");
	        $display ("To avoid this, please set PLLOUT_PHASE = \"NONE\" ");
	        $display ("******************************************************************");
		end
	end
 else
 		begin
	        $display ("************************SBT : Attention***************************");
	        $display ("Please set FEEDBACK_PATH to a valid value. Legal settings should be one of \"SIMPLE\", \"DELAY\", \"PHASE_AND_DELAY\", \"EXTERNAL\"");
	        $display ("******************************************************************");
  end 
end


mux4to1 instShftRegOutSelMux (
      .a (phase0net),
      .b (phase90net),
      .c (phase180net),
      .d (phase270net),
      .select (phasesel[1:0]),
      .o (phaseShiftMuxOutNet)
		);

ShiftReg instShftReg (
		.clk (ABPLLOUT),
		.init (RESET),
		.phase0 (phase0net),
		.phase90  (phase90net),
		.phase180 (phase180net),
		.phase270 (phase270net)
		);

mux4to1 instDlyAdjInMux (
		.a (ABPLLOUT),
		.b (phase0net),
		.c (phase0net),
		.d (EXTFEEDBACK),
		.select (delaymuxsel[1:0]),
		.o (finedelayin)
		);


FineDlyAdj instFineDlyAdj (
		.DlyAdj (DYNAMICDELAY),
		.signalin (finedelayin),
		.delayedout (finedelayout)
		);
defparam instFineDlyAdj.FIXED_DELAY_ADJUSTMENT = FIXED_DELAY_ADJUSTMENT;
defparam instFineDlyAdj.DELAY_ADJUSTMENT_MODE = DELAY_ADJUSTMENT_MODE;


 //buf #1750 (finedelayout, finedelayin);

ABIPTBS8 instABitsPLL (
		.REF (REFERENCECLK),
		.FB (FBnet),
		.FSE (FSEnet),
		.BYPASS (BYPASS),
		.RESET (RESET),
		.DIVF5 (DIVFBus[5]),
		.DIVF4 (DIVFBus[4]),
		.DIVF3 (DIVFBus[3]),
		.DIVF2 (DIVFBus[2]),
		.DIVF1 (DIVFBus[1]),
		.DIVF0 (DIVFBus[0]),
		.DIVQ2 (DIVQBus[2]),
		.DIVQ1 (DIVQBus[1]),
		.DIVQ0 (DIVQBus[0]),
		.DIVR3 (DIVRBus[3]),
		.DIVR2 (DIVRBus[2]),
		.DIVR1 (DIVRBus[1]),
		.DIVR0 (DIVRBus[0]),
		.RANGE2 (RANGEBus[2]),
		.RANGE1 (RANGEBus[1]),
		.RANGE0 (RANGEBus[0]),

		.LOCK (LOCK),
		.PLLOUT (ABPLLOUT)
		);

endmodule //SbtSPLL




`timescale 1ps/1ps
module SB_PLL_CORE (
		REFERENCECLK,		//Driven by core logic
		PLLOUTCORE,		//PLL output to core logic
		PLLOUTGLOBAL,	   	//PLL output to global network
		EXTFEEDBACK,  			//Driven by core logic
		DYNAMICDELAY,		//Driven by core logic
		LOCK,				//Output of PLL
		BYPASS,				//Driven by core logic
		RESET,				//Driven by core logic
		SDI,				//Driven by core logic. Test Pin
		SDO,				//Output to RB Logic Tile. Test Pin
		SCLK,				//Driven by core logic. Test Pin
		LATCHINPUTVALUE 	//iCEGate signal
);
input 	REFERENCECLK;		//Driven by core logic
output 	PLLOUTCORE;		//PLL output to core logic
output	PLLOUTGLOBAL;	   	//PLL output to global network
input	EXTFEEDBACK;  			//Driven by core logic
input	[3:0] DYNAMICDELAY;  	//Driven by core logic
output	LOCK;				//Output of PLL
input	BYPASS;				//Driven by core logic
input	RESET;				//Driven by core logic
input	LATCHINPUTVALUE; 	//iCEGate signal
//Test Pins
output	SDO;				//Output of PLL
input	SDI;				//Driven by core logic
input	SCLK;				//Driven by core logic

//Frequency Specification
//parameter REFERENCE_CLK_FREQUENCY = 100; 		//Floating Point
//parameter PLLOUT_FREQUENCY = 100;			//Floating Point
//parameter REFERENCE_CLK_DIVIDE_BY = 1;  		//Integer  Hide these for now
//parameter REFERENCE_CLK_MULTIPLY_BY = 1; 		//Integer  Hide these for now

//Feedback
parameter FEEDBACK_PATH = "SIMPLE";	//String  (simple, delay, phase_and_delay, external) (3 cbits, not 2)
parameter DELAY_ADJUSTMENT_MODE = "DYNAMIC"; 
parameter FIXED_DELAY_ADJUSTMENT = 0; 		//Integer. 
parameter PLLOUT_PHASE = "NONE"; //0deg,90deg,180deg,270deg,none

//Use the Spreadsheet to populate the values below.
parameter DIVR = 4'b0000; 	//determine a good default value
parameter DIVF = 6'b000000; //determine a good default value
parameter DIVQ = 3'b000; 	//determine a good default value
parameter FILTER_RANGE = 3'b000; 	//determine a good default value

//Additional cbits
parameter ENABLE_ICEGATE = 1'b0;

//Test Mode parameter
parameter TEST_MODE = 1'b0;
parameter EXTERNAL_DIVIDE_FACTOR = 1; //Not used by model. Added for PLL Config GUI.


SbtSPLL instSbtSPLL (
		.REFERENCECLK (REFERENCECLK),		//Driven by core logic
		.EXTFEEDBACK (EXTFEEDBACK),  			//Driven by core logic
		.DYNAMICDELAY (DYNAMICDELAY),		//Driven by core logic
		.BYPASS (BYPASS),				//Driven by core logic
		.RESET (~RESET),				//Driven by core logic
		
		.PLLOUT (SPLLOUTnet),		//PLL output to core logic
		.LOCK (LOCK)   		//Output of PLL

);
defparam instSbtSPLL.DIVR = DIVR;	
defparam instSbtSPLL.DIVF = DIVF;
defparam instSbtSPLL.DIVQ = DIVQ;
defparam instSbtSPLL.FILTER_RANGE = FILTER_RANGE;
defparam instSbtSPLL.FEEDBACK_PATH = FEEDBACK_PATH;
defparam instSbtSPLL.DELAY_ADJUSTMENT_MODE = DELAY_ADJUSTMENT_MODE;
defparam instSbtSPLL.FIXED_DELAY_ADJUSTMENT = FIXED_DELAY_ADJUSTMENT; 
defparam instSbtSPLL.PLLOUT_PHASE = PLLOUT_PHASE;


assign PLLOUTCORE = ((ENABLE_ICEGATE != 0) && LATCHINPUTVALUE) ? PLLOUTCORE : SPLLOUTnet;
assign PLLOUTGLOBAL = ((ENABLE_ICEGATE != 0) && LATCHINPUTVALUE)  ? PLLOUTGLOBAL : SPLLOUTnet;

`ifdef TIMINGCHECK
specify
   (REFERENCECLK *> PLLOUTGLOBAL) = (1.0, 1.0);
   (REFERENCECLK *> PLLOUTCORE) = (1.0, 1.0);
endspecify
`endif

endmodule // SB_PLL_CORE



`timescale 1ps/1ps
module SB_PLL_PAD (
		PACKAGEPIN,		//Driven by core logic
		PLLOUTCORE,		//PLL output to core logic
		PLLOUTGLOBAL,	   	//PLL output to global network
		EXTFEEDBACK,  			//Driven by core logic
		DYNAMICDELAY,		//Driven by core logic
		LOCK,				//Output of PLL
		BYPASS,				//Driven by core logic
		RESET,				//Driven by core logic
		SDI,				//Driven by core logic. Test Pin
		SDO,				//Output to RB Logic Tile. Test Pin
		SCLK,				//Driven by core logic. Test Pin
		LATCHINPUTVALUE 	//iCEGate signal
);
inout 	PACKAGEPIN;		//Driven by core logic
output 	PLLOUTCORE;		//PLL output to core logic
output	PLLOUTGLOBAL;	   	//PLL output to global network
input	EXTFEEDBACK;  			//Driven by core logic
input	[3:0] DYNAMICDELAY;  	//Driven by core logic
output	LOCK;				//Output of PLL
input	BYPASS;				//Driven by core logic
input	RESET;				//Driven by core logic
input	LATCHINPUTVALUE; 	//iCEGate signal
//Test Pins
output	SDO;				//Output of PLL
input	SDI;				//Driven by core logic
input	SCLK;				//Driven by core logic

//Frequency Specification
//parameter REFERENCE_CLK_FREQUENCY = 100; 		//Floating Point
//parameter PLLOUT_FREQUENCY = 100;			//Floating Point

//Feedback
parameter FEEDBACK_PATH = "SIMPLE";	//String  (simple, delay, phase_and_delay, external) (3 cbits, not 2)
parameter DELAY_ADJUSTMENT_MODE = "DYNAMIC"; //String. 
parameter FIXED_DELAY_ADJUSTMENT = 0; 		//Integer. 
parameter PLLOUT_PHASE = "NONE"; //0deg,90deg,180deg,270deg,none

//Use the Spreadsheet to populate the values below.
parameter DIVR = 4'b0000; 	//determine a good default value
parameter DIVF = 6'b000000; //determine a good default value
parameter DIVQ = 3'b000; 	//determine a good default value
parameter FILTER_RANGE = 3'b000; 	//determine a good default value

//Additional cbits
parameter ENABLE_ICEGATE = 1'b0;

//Test Mode parameter
parameter TEST_MODE = 1'b0;
parameter EXTERNAL_DIVIDE_FACTOR = 1; //Not used by model. Added for PLL Config GUI.

SbtSPLL instSbtSPLL (
		.REFERENCECLK (PACKAGEPIN),		//Driven by core logic
		.EXTFEEDBACK (EXTFEEDBACK),  			//Driven by core logic
		.DYNAMICDELAY (DYNAMICDELAY),		//Driven by core logic
		.BYPASS (BYPASS),				//Driven by core logic
		.RESET (~RESET),				//Driven by core logic
		
		.PLLOUT (SPLLOUTnet),		//PLL output to core logic
		.LOCK (LOCK)   		//Output of PLL
);
defparam instSbtSPLL.DIVR = DIVR;	
defparam instSbtSPLL.DIVF = DIVF;
defparam instSbtSPLL.DIVQ = DIVQ;
defparam instSbtSPLL.FILTER_RANGE = FILTER_RANGE;
defparam instSbtSPLL.FEEDBACK_PATH = FEEDBACK_PATH;
defparam instSbtSPLL.DELAY_ADJUSTMENT_MODE = DELAY_ADJUSTMENT_MODE;
defparam instSbtSPLL.FIXED_DELAY_ADJUSTMENT = FIXED_DELAY_ADJUSTMENT; 
defparam instSbtSPLL.PLLOUT_PHASE = PLLOUT_PHASE;


assign PLLOUTCORE = ((ENABLE_ICEGATE != 0) && LATCHINPUTVALUE) ? PLLOUTCORE : SPLLOUTnet;
assign PLLOUTGLOBAL = ((ENABLE_ICEGATE != 0) && LATCHINPUTVALUE)  ? PLLOUTGLOBAL : SPLLOUTnet;

`ifdef TIMINGCHECK
specify
   (PACKAGEPIN *> PLLOUTGLOBAL) = (1.0, 1.0);
   (PACKAGEPIN *> PLLOUTCORE) = (1.0, 1.0);

endspecify
`endif

endmodule // SB_PLL_PAD



`timescale 1ps/1ps
module SB_PLL_2_PAD (
		PACKAGEPIN,		//Driven by core logic
		PLLOUTCOREA,		//DIN0 output to core logic
		PLLOUTGLOBALA,	   	//GLOBALOUTPUTBUFFER
        PLLOUTCOREB,		//PLL output to core logic
		PLLOUTGLOBALB,	   	//PLL output to global network
		EXTFEEDBACK,  			//Driven by core logic
		DYNAMICDELAY,		//Driven by core logic
		LOCK,				//Output of PLL
		BYPASS,				//Driven by core logic
		RESET,				//Driven by core logic
		SDI,				//Driven by core logic. Test Pin
		SDO,				//Output to RB Logic Tile. Test Pin
		SCLK,				//Driven by core logic. Test Pin
		LATCHINPUTVALUE 	//iCEGate signal
);
inout 	PACKAGEPIN;		//Driven by core logic
output  PLLOUTCOREA;		//PLL output to core logic
output	PLLOUTGLOBALA;	   	//PLL output to global network
output  PLLOUTCOREB;		//PLL output to core logic
output	PLLOUTGLOBALB;	   	//PLL output to global network
input	EXTFEEDBACK;  			//Driven by core logic
input	[3:0] DYNAMICDELAY;  	//Driven by core logic
output	LOCK;				//Output of PLL
input	BYPASS;				//Driven by core logic
input	RESET;				//Driven by core logic
input	LATCHINPUTVALUE; 	//iCEGate signal
//Test Pins
output	SDO;				//Output of PLL
input	SDI;				//Driven by core logic
input	SCLK;				//Driven by core logic

//Frequency Specification
//parameter REFERENCE_CLK_FREQUENCY = 100; 		//Floating Point
//parameter PLLOUT_FREQUENCY_PORTB = 100;			//Floating Point

//Feedback
parameter FEEDBACK_PATH = "SIMPLE";	//simple, delay, phase_and_delay, external 
parameter DELAY_ADJUSTMENT_MODE = "DYNAMIC"; //Fixed, Dynamic 
parameter FIXED_DELAY_ADJUSTMENT = 0; 		// 0-15 
parameter PLLOUT_PHASE = "NONE"; //0deg,90deg,180deg,270deg,none

//Use the Spreadsheet to populate the values below.
parameter DIVR = 4'b0000; 	//determine a good default value
parameter DIVF = 6'b000000; //determine a good default value
parameter DIVQ = 3'b000; 	//determine a good default value
parameter FILTER_RANGE = 3'b000; 	//determine a good default value

//Additional cbits
parameter ENABLE_ICEGATE_PORTA = 1'b0;
parameter ENABLE_ICEGATE_PORTB = 1'b0;

//Test Mode parameter
parameter TEST_MODE = 1'b0;
parameter EXTERNAL_DIVIDE_FACTOR = 1; //Not used by model. Added for PLL Config GUI.

SbtSPLL instSbtSPLL (
		.REFERENCECLK (PACKAGEPIN),		//Driven by core logic
		.EXTFEEDBACK (EXTFEEDBACK),  			//Driven by core logic
		.DYNAMICDELAY (DYNAMICDELAY),		//Driven by core logic
		.BYPASS (BYPASS),				//Driven by core logic
		.RESET (~RESET),				//Driven by core logic
		
		.PLLOUT (SPLLOUTnet),		//PLL output to core logic
		.LOCK (LOCK)   		//Output of PLL
);
defparam instSbtSPLL.DIVR = DIVR;	
defparam instSbtSPLL.DIVF = DIVF;
defparam instSbtSPLL.DIVQ = DIVQ;
defparam instSbtSPLL.FILTER_RANGE = FILTER_RANGE;
defparam instSbtSPLL.FEEDBACK_PATH = FEEDBACK_PATH;
defparam instSbtSPLL.DELAY_ADJUSTMENT_MODE = DELAY_ADJUSTMENT_MODE;
defparam instSbtSPLL.FIXED_DELAY_ADJUSTMENT = FIXED_DELAY_ADJUSTMENT; 
defparam instSbtSPLL.PLLOUT_PHASE = PLLOUT_PHASE;


assign PLLOUTCOREA = ((ENABLE_ICEGATE_PORTA != 0) && LATCHINPUTVALUE) ? PLLOUTCOREA : PACKAGEPIN;
assign PLLOUTGLOBALA = ((ENABLE_ICEGATE_PORTA != 0) && LATCHINPUTVALUE)  ? PLLOUTGLOBALA : PACKAGEPIN;
assign PLLOUTCOREB = ((ENABLE_ICEGATE_PORTB != 0) && LATCHINPUTVALUE) ? PLLOUTCOREB : SPLLOUTnet;
assign PLLOUTGLOBALB = ((ENABLE_ICEGATE_PORTB != 0) && LATCHINPUTVALUE)  ? PLLOUTGLOBALB : SPLLOUTnet;

`ifdef TIMINGCHECK
specify
   (PACKAGEPIN *> PLLOUTGLOBALA) = (1.0, 1.0);
   (PACKAGEPIN *> PLLOUTCOREA) = (1.0, 1.0);
   (PACKAGEPIN *> PLLOUTGLOBALB) = (1.0, 1.0);
   (PACKAGEPIN *> PLLOUTCOREB) = (1.0, 1.0);

endspecify
`endif

endmodule // SB_PLL_2_PAD



/****** ice40 PLL prims*****/
////////////////////////////////////////////////////////
/////		Static PLL Model 	////////////////
////////////////////////////////////////////////////////
/*

`timescale 1ps/1ps

module ShiftReg427 (clk, init, phase0, phase90);
input clk, init; 
output phase0, phase90;

parameter SHIFTREG_DIV_MODE = 2'b00; // 00-->Divide by 4 ,  01-->Divide by 7 , 
				     //	10 --> "INVALID mode" , 11--> Divide by 5(HDMI).
//parameter SHIFTREG_DIV_MODE = 1'b0; //0-->Divide by 4, 1-->Divide by 7.

reg ff1, ff2, ff3, ff4, ff5, ff6, ff7;

always @ (posedge clk or posedge init)
   begin
	if (init)  
		begin
			ff1	 = 1'b0;
			ff2	 = 1'b0;
			ff3	 = 1'b0;
			ff4	 = 1'b1;
			ff5	 = 1'b1;
			ff6	 = 1'b1;
			ff7	 = 1'b1;
		end
	else	
		begin
	   	    	ff1 <= ff7;
			ff2 <= ff1;
			ff3 <= ff2;
			ff4 <= ff3;
		//	ff5 <= ff4;
			if 	(SHIFTREG_DIV_MODE == 2'b00)
			begin 
				ff5 <= ff4; 
				ff6 <= ff2;
			end 
			else if (SHIFTREG_DIV_MODE == 2'b01)
			begin 
				ff5 <= ff4; 
				ff6 <= ff5;
			end 
			else if (SHIFTREG_DIV_MODE == 2'b11)
			begin
				ff5 <= ff2; 
				ff6 <= ff5;
			end 
			else if (SHIFTREG_DIV_MODE == 2'b10) 
			begin 
				$display("Incorrect SHIFTREG_DIV_MODE set for simulation\n");
				$finish; 
			end 

			ff7 <= ff6;
		end
    end

assign phase0 = ff1;
assign phase90 = ff2;

endmodule
*/

/*
`timescale 1ps/1ps
module SbtSPLL40 (
		REFERENCECLK,
		EXTFEEDBACK,
		DYNAMICDELAY,
		BYPASS,	
		RESETB,		
		
		PLLOUT1,		
		PLLOUT2,		
		LOCK   		
);

//----------------------------------------------------------------------
// Port Declarations
//----------------------------------------------------------------------

// Inputs

input REFERENCECLK;		
input	EXTFEEDBACK;  
input	[7:0] DYNAMICDELAY;  
input	BYPASS;				
input	RESETB;			

// Outputs
output 	PLLOUT1, PLLOUT2;	
output	LOCK;				//Output of PLL

//Feedback
parameter FEEDBACK_PATH = "SIMPLE";	//String  (simple, delay, phase_and_delay, external) 
parameter DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED"; 
parameter DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED"; 
parameter SHIFTREG_DIV_MODE = 2'b00; //00-->Divide by 4, 01-->Divide by 7 , 10 --> invalid , 11 --> Divide by 5 (HDMI).
//parameter SHIFTREG_DIV_MODE = 1'b0; //0-->Divide by 4, 1-->Divide by 7.
parameter FDA_FEEDBACK = 4'b0000; 		//Integer. 

//Output 
parameter FDA_RELATIVE = 4'b0000; 		//Integer. 
parameter PLLOUT_SELECT_PORTA = "GENCLK"; //
parameter PLLOUT_SELECT_PORTB = "GENCLK"; //

//Use the Spreadsheet to populate the values below.
parameter DIVR = 4'b0000; 	//determine a good default value
parameter DIVF = 7'b0000000; //determine a good default value
parameter DIVQ = 3'b000; 	//determine a good default value
parameter FILTER_RANGE = 3'b000; 	//determine a good default value

//Additional cbits
parameter ENBLE_ICEGATE_PORTA = 1'b0;
parameter ENABLE_ICEGATE_PORTB = 1'b0;


wire FSEnet;
wire FBnet;
wire finedelayFBin, finedelayFBout;
//wire [5:0] DIVFBus = DIVF; 
wire [6:0] DIVFBus = DIVF; 
wire [3:0] DIVRBus = DIVR; 
wire [2:0] DIVQBus = DIVQ; 
wire [2:0] RANGEBus = FILTER_RANGE; 
wire ABPLLOUT;
reg [1:0] pllout1Sel;
reg [1:0] pllout2Sel;
reg [1:0] delaymuxsel;
reg ABPLLOUTDiv2;

//reg fbout;

initial
begin
  ABPLLOUTDiv2 = 1'b0;
end

always @ (posedge ABPLLOUT)
	ABPLLOUTDiv2 = ~ABPLLOUTDiv2;


initial
begin
 if (PLLOUT_SELECT_PORTA == "SHIFTREG_0deg")
    pllout1Sel = 2'b00;
else if (PLLOUT_SELECT_PORTA == "SHIFTREG_90deg")
    pllout1Sel = 2'b01;
else if (PLLOUT_SELECT_PORTA == "GENCLK_HALF")
    pllout1Sel = 2'b10;
else if (PLLOUT_SELECT_PORTA == "GENCLK")
    pllout1Sel = 2'b11;
else 
   begin
	        $display ("************************SBT : ERROR ****************************");
	        $display ("Parameter PLLOUT_SELECT_PORTA is set to an illegal value.");
	        $display ("Legal values should be one of \"SHIFTREG_0deg\", \"SHIFTREG_90deg\", \"GENCLK_HALF\", \"GENCLK\". ");
	        $display ("Due to incorrect configuration of the PLL, the simulation results are invalid.");
	        $display ("****************************************************************");
	        $finish;
   end
end

initial
begin
 if (PLLOUT_SELECT_PORTB == "SHIFTREG_0deg")
    pllout2Sel = 2'b00;
else if (PLLOUT_SELECT_PORTB == "SHIFTREG_90deg")
    pllout2Sel = 2'b01;
else if (PLLOUT_SELECT_PORTB == "GENCLK_HALF")
    pllout2Sel = 2'b10;
else if (PLLOUT_SELECT_PORTB == "GENCLK")
    pllout2Sel = 2'b11;
else 
   begin
	        $display ("************************SBT : ERROR ****************************");
	        $display ("Parameter PLLOUT_SELECT_PORTB is set to an illegal value.");
	        $display ("Legal values should be one of \"SHIFTREG_0deg\", \"SHIFTREG_90deg\", \"GENCLK_HALF\", \"GENCLK\". ");
	        $display ("Due to incorrect configuration of the PLL, the simulation results are invalid.");
	        $display ("****************************************************************");
	        $finish;
   end
end

assign FSEnet = (FEEDBACK_PATH == "SIMPLE") ? 1'b1 : 1'b0;
assign FBnet = (FEEDBACK_PATH == "SIMPLE") ? 1'b0 : finedelayFBout;


initial
begin

 if (FEEDBACK_PATH != "EXTERNAL")
 	begin
	    $display ("************************SBT : Info*****************************");
	    $display ("Note that any signal connection to the EXTFEEDBACK port of the PLL will be ignored");
	    $display ("***************************************************************");
	   	end
 if (FEEDBACK_PATH == "EXTERNAL")
    begin 
       delaymuxsel = 2'b11;
        if ( (DELAY_ADJUSTMENT_MODE_FEEDBACK != "FIXED") && (DELAY_ADJUSTMENT_MODE_FEEDBACK != "DYNAMIC") )
		begin
	        $display ("************************SBT : ERROR ************************");
	        $display ("Since FEEDBACK_PATH=\"EXTERNAL\", DELAY_ADJUSTMENT_MODE_FEEDBACK should be \"FIXED\" or \"DYNAMIC\"");
	        $display ("Due to incorrect configuration of the PLL, the simulation results are invalid.");
	        $display ("***************************************************************");
	        $finish;
		end
		if (PLLOUT_SELECT_PORTA == "SHIFTREG_0deg" || PLLOUT_SELECT_PORTA == "SHIFTREG_90deg"
		    || PLLOUT_SELECT_PORTB == "SHIFTREG_0deg" || PLLOUT_SELECT_PORTB == "SHIFTREG_90deg")  // model divby2 clk, check changed params, compile
		begin
	        $display ("************************ SBT : ERROR **************************");
	        $display ("Since FEEDBACK_PATH=\"EXTERNAL\", Phase Adjustment is NOT permitted.");
	        $display ("*************************************************************");
	        $finish;
		end
    end				
 else if (FEEDBACK_PATH == "DELAY")
    begin 
    	delaymuxsel = 2'b00;
        if ( (DELAY_ADJUSTMENT_MODE_FEEDBACK != "FIXED") && (DELAY_ADJUSTMENT_MODE_FEEDBACK != "DYNAMIC") )
		begin
	        $display ("************************ SBT : ERROR **************************");
	        $display ("Since FEEDBACK_PATH=\"DELAY\", DELAY_ADJUSTMENT_MODE_FEEDBACK should be \"FIXED\" or \"DYNAMIC\"");
	        $display ("Due to incorrect configuration of the PLL, the simulation results are invalid.");
	        $display ("***************************************************************");
	        $finish;
		end
		if (PLLOUT_SELECT_PORTA == "SHIFTREG_0deg" || PLLOUT_SELECT_PORTA == "SHIFTREG_90deg"
		    || PLLOUT_SELECT_PORTB == "SHIFTREG_0deg" || PLLOUT_SELECT_PORTB == "SHIFTREG_90deg")  //use PLLOUT_SELECT, model divby2 clk, check changed params, compile
		begin
	        $display ("************************ SBT : ERROR **************************");
	        $display ("Since FEEDBACK_PATH=\"DELAY\", Phase Adjustment is NOT permitted. Please set PLLOUT_SELECT_PORTA/B=\"GENCLK\" or \"GENCLK_HALF\"");
		    $display ("Due to incorrect configuration of the PLL, the simulation results are invalid.");
	        $display ("***************************************************************");
	        $finish;
		end
    end				
 else if (FEEDBACK_PATH == "PHASE_AND_DELAY")
	begin
    	delaymuxsel = 2'b01;
        if ( (DELAY_ADJUSTMENT_MODE_FEEDBACK != "FIXED") && (DELAY_ADJUSTMENT_MODE_FEEDBACK != "DYNAMIC") )
		begin
	        $display ("************************SBT : Attention************************");
	        $display ("Since FEEDBACK_PATH=\"PHASE_AND_DELAY\", DELAY_ADJUSTMENT_MODE_FEEDBACK should be FIXED or DYNAMIC");
	        $display ("***************************************************************");
		end
		if ( (PLLOUT_SELECT_PORTA != "SHIFTREG_0deg") && (PLLOUT_SELECT_PORTA != "SHIFTREG_90deg" )
				&& (PLLOUT_SELECT_PORTB != "SHIFTREG_0deg") && (PLLOUT_SELECT_PORTB != "SHIFTREG_90deg") )
		begin
	        $display ("************************SBT : Attention************************");
	        $display ("FEEDBACK_PATH=\"PHASE_AND_DELAY\", but PLLOUT_SELECT_PORTA/B is not specified correctly");
	        $display ("***************************************************************");
		end
    end				
else if (FEEDBACK_PATH == "SIMPLE")
   begin
		//Ignore DELAY_ADJUSTMENT_MODE_FEEDBACK, FDA_FEEDBACK   
	  $display ("************************SBT : Attention***************************");
	  $display ("Since FEEDBACK_PATH=\"SIMPLE\", the FDA_FEEDBACK value will be ignored");
	  $display ("******************************************************************");


	if (PLLOUT_SELECT_PORTA == "SHIFTREG_0deg" || PLLOUT_SELECT_PORTA == "SHIFTREG_90deg"
		    || PLLOUT_SELECT_PORTB == "SHIFTREG_0deg" || PLLOUT_SELECT_PORTB == "SHIFTREG_90deg")  //use PLLOUT_SELECT, model divby2 clk, check changed params, compile
		begin
	        $display ("************************SBT : Attention***************************");
	        $display ("The PLL output frequency will be divided by 4 or 7 and phase shifted.");
	        $display ("To avoid this, please set PLLOUT_SELECT_PORTA/B = \"GENCLK\" ");
	        $display ("******************************************************************");
		end
	end
 else
 		begin
	        $display ("************************SBT : Attention***************************");
	        $display ("Please set FEEDBACK_PATH to a valid value. Legal settings should be one of \"SIMPLE\", \"DELAY\", \"PHASE_AND_DELAY\", \"EXTERNAL\"");
	        $display ("******************************************************************");
  end 

	if( SHIFTREG_DIV_MODE == 2'b10) 
		begin
	        $display ("************************ SBT : ERROR **************************");
	        $display ("SHIFTREG_DIV_MODE = 2'b10 is NOT permitted. Please set it 2'b00/2'b01/2'b11");
	        $display ("Due to incorrect configuration of the PLL, the simulation results are invalid.");
	        $display ("***************************************************************");
	        $finish;
		end 
   	
end


ShiftReg427 instShftReg427 (
		.clk (ABPLLOUT),
		.init (RESETB),
		.phase0 (phase0net),
		.phase90 (phase90net)
		);
defparam instShftReg427.SHIFTREG_DIV_MODE = SHIFTREG_DIV_MODE;

mux4to1 instFBDlyAdjInMux (
		.a (ABPLLOUT),
		.b (phase0net),
		.c (phase0net),
		.d (EXTFEEDBACK),
		.select (delaymuxsel[1:0]),
		.o (finedelayFBin)
		);


mux4to1 instPLLOUT2SelMux (
		.a (phase0net),
		.b (phase90net),
		.d(ABPLLOUT),
		.c (ABPLLOUTDiv2),
		.select (pllout2Sel[1:0]),
		.o (pllout2Muxnet)
		);
assign PLLOUT2 = (BYPASS == 1'b1) ? REFERENCECLK : pllout2Muxnet;

mux4to1 instPLLOUT1SelMux (
		.a (phase0net),
		.b (phase90net),
		.d (ABPLLOUT),
		.c (ABPLLOUTDiv2),
		.select (pllout1Sel[1:0]),
		.o (pllout1Muxnet)
		);
assign fdaRelInput = (BYPASS == 1'b1) ? REFERENCECLK : pllout1Muxnet;


FineDlyAdj instFineDlyAdjFB (
		.DlyAdj (DYNAMICDELAY[3:0]),
		.signalin (finedelayFBin),
		.delayedout (finedelayFBout)
		);
defparam instFineDlyAdjFB.FIXED_DELAY_ADJUSTMENT = FDA_FEEDBACK;
defparam instFineDlyAdjFB.DELAY_ADJUSTMENT_MODE = DELAY_ADJUSTMENT_MODE_FEEDBACK;

FineDlyAdj instFineDlyAdjRel (
		.DlyAdj (DYNAMICDELAY[7:4]),
		.signalin (fdaRelInput),
		.delayedout (PLLOUT1)
		);
defparam instFineDlyAdjRel.FIXED_DELAY_ADJUSTMENT = FDA_RELATIVE;
defparam instFineDlyAdjRel.DELAY_ADJUSTMENT_MODE = DELAY_ADJUSTMENT_MODE_RELATIVE;


ABIWTCZ4 instABitsPLL (
		.REF (REFERENCECLK),
		.FB (FBnet),
		.FSE (FSEnet),
		.BYPASS (BYPASS),
		.RESET (RESETB),
		.DIVF6 (DIVFBus[6]),
		.DIVF5 (DIVFBus[5]),
		.DIVF4 (DIVFBus[4]),
		.DIVF3 (DIVFBus[3]),
		.DIVF2 (DIVFBus[2]),
		.DIVF1 (DIVFBus[1]),
		.DIVF0 (DIVFBus[0]),
		.DIVQ2 (DIVQBus[2]),
		.DIVQ1 (DIVQBus[1]),
		.DIVQ0 (DIVQBus[0]),
		.DIVR3 (DIVRBus[3]),
		.DIVR2 (DIVRBus[2]),
		.DIVR1 (DIVRBus[1]),
		.DIVR0 (DIVRBus[0]),
		.RANGE2 (RANGEBus[2]),
		.RANGE1 (RANGEBus[1]),
		.RANGE0 (RANGEBus[0]),

		.LOCK (LOCK),
		.PLLOUT (ABPLLOUT)
		);

endmodule //SbtSPLL
*/ 


////////////////////////////////////////////////////////
/////		Dynamic PLL Model 	////////////////
////////////////////////////////////////////////////////
/* 
`timescale 1ps/1ps
module pllcfg_dynamicsetting_shiftreg (pll_sck,pll_sdi, q);
input pll_sck, pll_sdi; 
output [26:0] q;

reg [26:0] q = 27'b0;

always @ (negedge pll_sck)
   begin
	 q[26:0] <= {q[25:0],pll_sdi};
   end

endmodule


`timescale 1ps/1ps 
module ShiftReg427_DS (clk, init, phase0, phase90, shiftregister_div_mode_sel);
input clk, init; 

output phase0, phase90;

//// parameter SHIFTREG_DIV_MODE = 2'b00; 
////					 00--> Divide by 4,
////					 01--> Divide by 7, 
//// 			     		 10--> INVALID mode, 
////					 11--> Divide by 5(HDMI).

input [1:0] shiftregister_div_mode_sel;

reg ff1, ff2, ff3, ff4, ff5, ff6, ff7;

always @ (posedge clk or posedge init)
   begin
	if (init)  
		begin
			ff1	 = 1'b0;
			ff2	 = 1'b0;
			ff3	 = 1'b0;
			ff4	 = 1'b1;
			ff5	 = 1'b1;
			ff6	 = 1'b1;
			ff7	 = 1'b1;
		end
	else	
		begin
	   	    	ff1 <= ff7;
			ff2 <= ff1;
			ff3 <= ff2;
			ff4 <= ff3;
		//	ff5 <= ff4;
			if 	(shiftregister_div_mode_sel == 2'b00)
			begin 
				ff5 <= ff4; 
				ff6 <= ff2;
			end 
			else if (shiftregister_div_mode_sel == 2'b01)
			begin 
				ff5 <= ff4; 
				ff6 <= ff5;
			end 
			else if (shiftregister_div_mode_sel == 2'b11)
			begin
				ff5 <= ff2; 
				ff6 <= ff5;
			end 
			else if (shiftregister_div_mode_sel == 2'b10) 
			begin 
				$display("Incorrect SHIFTREG_DIV_MODE set for simulation\n");
				$finish; 
			end 

			ff7 <= ff6;
		end
    end

assign phase0 = ff1;
assign phase90 = ff2;

endmodule

//Sbt Dynamic Setting PLL40 
module Sbt_DS_PLL40 (
		PACKAGEPIN,		//Driven by IO clock
		CORE_REF_CLK,		//Driven by core logic
		EXTFEEDBACK,
		DYNAMICDELAY,
		BYPASS,	
		RESETB,		
		
		PLL_SCK,
		PLL_SDI,
		PLL_SDO,
		
		PLLOUT1,		
		PLLOUT2,		
		LOCK   		
);

//----------------------------------------------------------------------
// Port Declarations
//----------------------------------------------------------------------
// Inputs
input 	PACKAGEPIN;			//Driven by IO clock
input 	CORE_REF_CLK;			//Driven by core logic
input	EXTFEEDBACK;  
input	[7:0] DYNAMICDELAY;  
input	BYPASS;				
input	RESETB;			
input	PLL_SCK;			
input	PLL_SDI;			

// Outputs
output 	PLLOUT1, PLLOUT2;	
output	LOCK;				
output	PLL_SDO;			

//----------------------------------------------------------------------
// ALL the parameter definitions here are just for STA timing analysis presume user will use those settings in the shift registers
//----------------------------------------------------------------------
//Feedback
parameter FEEDBACK_PATH = "SIMPLE";			//String  (simple, delay, phase_and_delay, external) 
parameter DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED"; 
parameter DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED"; 
parameter SHIFTREG_DIV_MODE = 2'b00; 			//00-->Divide by 4, 01-->Divide by 7 , 10 --> invalid , 11 --> Divide by 5 (HDMI).
//parameter SHIFTREG_DIV_MODE = 1'b0; 			//0-->Divide by 4, 1-->Divide by 7.
parameter FDA_FEEDBACK = 4'b0000; 			//Integer. 

//Output 
parameter FDA_RELATIVE = 4'b0000; 			//Integer. 
parameter PLLOUT_SELECT_PORTA = "GENCLK"; 		
parameter PLLOUT_SELECT_PORTB = "GENCLK";		
//Use the Spreadsheet to populate the values below.
parameter DIVR = 4'b0000; 				//determine a good default value
parameter DIVF = 7'b0000000; 				//determine a good default value
parameter DIVQ = 3'b000; 				//determine a good default value
parameter FILTER_RANGE = 3'b000; 			//determine a good default value

//Additional cbits
parameter ENBLE_ICEGATE_PORTA = 1'b0;
parameter ENABLE_ICEGATE_PORTB = 1'b0;


parameter TEST_MODE = 1'b1;				//TEST_MODE has to be set to "1" for PLL dynamic setting

wire  [26:0] PLLCFG_SREG;
wire FSEnet = PLLCFG_SREG[25];
wire FBnet;
wire finedelayFBin, finedelayFBout;
// change for shift register dynamic PLL setting 
wire [6:0] DIVFBus = PLLCFG_SREG[10:4];			//DIVF; 
wire [3:0] DIVRBus = PLLCFG_SREG[3:0];			//DIVR; 
wire [2:0] DIVQBus = PLLCFG_SREG[13:11];		//DIVQ; 
wire [2:0] RANGEBus = PLLCFG_SREG[16:14];		//FILTER_RANGE; 
wire ABPLLOUT;
wire [1:0] pllout1Sel = PLLCFG_SREG[24:23];
wire [1:0] pllout2Sel = PLLCFG_SREG[20:19];
wire [1:0] shiftregister_div_mode_sel;			//SHIFTREG_DIV_MODE
// change for shift register dynamic PLL setting 
wire [1:0] delaymuxsel = PLLCFG_SREG[18:17];
reg ABPLLOUTDiv2;
wire REFERENCECLK;		

assign shiftregister_div_mode_sel =	{PLLCFG_SREG[26],PLLCFG_SREG[21]};	
assign FBnet = (FSEnet) ? 1'b0 : finedelayFBout;
assign PLL_SDO = PLLCFG_SREG[26];
assign REFERENCECLK = (PLLCFG_SREG[22]) ? CORE_REF_CLK : PACKAGEPIN;
//reg fbout;

reg [4:0] DS_POSCLK_COUNTER, DS_NEGCLK_COUNTER;
wire DS_NEGCLK_COUNTER_CLEAR;

initial
begin
	DS_POSCLK_COUNTER <=5'd27;
	DS_NEGCLK_COUNTER <=5'd27;
end

always @(negedge RESETB) 
begin
	DS_POSCLK_COUNTER <=5'd27;
	DS_NEGCLK_COUNTER <=5'd27;
end

always @(posedge PLL_SCK) 
begin
	if (DS_POSCLK_COUNTER == 5'b0)
	begin
        $display ("************************SBT : PLL_DS ERROR ****************************");
        $display ("Once the 27 cycles are completed, SCLK needs to stop.");
        $display ("****************************************************************");
        $finish;
	end
	else DS_POSCLK_COUNTER <= DS_POSCLK_COUNTER - 5'd1;
end

always @(negedge PLL_SCK) 
begin
	if (DS_NEGCLK_COUNTER == 5'b0)
	begin
        $display ("************************SBT : PLL_DS ERROR ****************************");
        $display ("Once the 27 cycles are completed, SCLK needs to stop.");
        $display ("****************************************************************");
        $finish;
	end
	else DS_NEGCLK_COUNTER <= DS_NEGCLK_COUNTER - 5'd1;
end

assign DS_NEGCLK_COUNTER_CLEAR = (DS_NEGCLK_COUNTER[4:0] == 5'b0);

always @(posedge PLL_SCK or negedge PLL_SCK) 
	if (RESETB == 0)
	begin
        $display ("************************SBT : PLL_DS ERROR ****************************");
        $display ("PLL RESETB needs to be held low while the data is shifted into the register by PLL_SCK clock.");
        $display ("****************************************************************");
        $finish;
	end

always @(posedge RESETB) 
	if ((DS_POSCLK_COUNTER != 5'b0) | (DS_NEGCLK_COUNTER != 5'b0))
	begin
        $display ("************************SBT : PLL_DS ERROR ****************************");
        $display ("Exactly 27 full clock cycles are needed to shift SDI data into the register.");
        $display ("****************************************************************");
        $finish;
	end

always @(posedge DS_NEGCLK_COUNTER_CLEAR) 
	begin
		# 10;
		if (RESETB == 1)
		begin
			$display ("************************SBT : PLL_DS ERROR ****************************");
			$display ("Release RESETB greater than 10ns once SCLK is stopped.");
			$display ("****************************************************************");
			$finish;
		end
	end

	
initial
begin
  ABPLLOUTDiv2 = 1'b0;
end

always @ (posedge ABPLLOUT)
	ABPLLOUTDiv2 = ~ABPLLOUTDiv2;


pllcfg_dynamicsetting_shiftreg instPLLCFG_DS_SReg(
		.pll_sck(PLL_SCK),
		.pll_sdi(PLL_SDI), 
		.q(PLLCFG_SREG)
		);

//shiftregister_div_mode_sel
//00-->Divide by 4, 01-->Divide by 7 , 10 --> invalid , 11 --> Divide by 5 (HDMI).
ShiftReg427_DS instShftReg427 (
		.clk (ABPLLOUT),
		.init (RESETB),
		.phase0 (phase0net),
		.phase90 (phase90net),
		.shiftregister_div_mode_sel(shiftregister_div_mode_sel)
		);

mux4to1 instFBDlyAdjInMux (
		.a (ABPLLOUT),
		.b (phase0net),
		.c (phase0net),
		.d (EXTFEEDBACK),
		.select (delaymuxsel[1:0]),
		.o (finedelayFBin)
		);


mux4to1 instPLLOUT2SelMux (
		.a (phase0net),
		.b (phase90net),
		.d(ABPLLOUT),
		.c (ABPLLOUTDiv2),
		.select (pllout2Sel[1:0]),
		.o (pllout2Muxnet)
		);
assign PLLOUT2 = (BYPASS == 1'b1) ? REFERENCECLK : pllout2Muxnet;

mux4to1 instPLLOUT1SelMux (
		.a (phase0net),
		.b (phase90net),
		.d (ABPLLOUT),
		.c (ABPLLOUTDiv2),
		.select (pllout1Sel[1:0]),
		.o (pllout1Muxnet)
		);
assign fdaRelInput = (BYPASS == 1'b1) ? REFERENCECLK : pllout1Muxnet;


FineDlyAdj instFineDlyAdjFB (
		.DlyAdj (DYNAMICDELAY[3:0]),
		.signalin (finedelayFBin),
		.delayedout (finedelayFBout)
		);
defparam instFineDlyAdjFB.FIXED_DELAY_ADJUSTMENT = FDA_FEEDBACK;
defparam instFineDlyAdjFB.DELAY_ADJUSTMENT_MODE = DELAY_ADJUSTMENT_MODE_FEEDBACK;

FineDlyAdj instFineDlyAdjRel (
		.DlyAdj (DYNAMICDELAY[7:4]),
		.signalin (fdaRelInput),
		.delayedout (PLLOUT1)
		);
defparam instFineDlyAdjRel.FIXED_DELAY_ADJUSTMENT = FDA_RELATIVE;
defparam instFineDlyAdjRel.DELAY_ADJUSTMENT_MODE = DELAY_ADJUSTMENT_MODE_RELATIVE;


ABIWTCZ4 instABitsPLL (
		.REF (REFERENCECLK),
		.FB (FBnet),
		.FSE (FSEnet),
		.BYPASS (BYPASS),
		.RESET (RESETB),
		.DIVF6 (DIVFBus[6]),
		.DIVF5 (DIVFBus[5]),
		.DIVF4 (DIVFBus[4]),
		.DIVF3 (DIVFBus[3]),
		.DIVF2 (DIVFBus[2]),
		.DIVF1 (DIVFBus[1]),
		.DIVF0 (DIVFBus[0]),
		.DIVQ2 (DIVQBus[2]),
		.DIVQ1 (DIVQBus[1]),
		.DIVQ0 (DIVQBus[0]),
		.DIVR3 (DIVRBus[3]),
		.DIVR2 (DIVRBus[2]),
		.DIVR1 (DIVRBus[1]),
		.DIVR0 (DIVRBus[0]),
		.RANGE2 (RANGEBus[2]),
		.RANGE1 (RANGEBus[1]),
		.RANGE0 (RANGEBus[0]),

		.LOCK (LOCK),
		.PLLOUT (ABPLLOUT)
		);

endmodule //Sbt_DS_PLL
*/ 


////-----------------------------------------------------
//// ------------ SB_PLL40_CORE  ------------------------
////-----------------------------------------------------

`timescale 1ps/1ps
module SB_PLL40_CORE (
		REFERENCECLK,			//Driven by core logic
		PLLOUTCORE,			//PLL output to core logic
		PLLOUTGLOBAL,	   		//PLL output to global network
		EXTFEEDBACK,  			//Driven by core logic
		DYNAMICDELAY,			//Driven by core logic
		LOCK,				//Output of PLL
		BYPASS,				//Driven by core logic
		RESETB,				//Driven by core logic
		SDI,				//Driven by core logic. Test Pin
		SDO,				//Output to RB Logic Tile. Test Pin
		SCLK,				//Driven by core logic. Test Pin
		LATCHINPUTVALUE 		//iCEGate signal
);

input 	REFERENCECLK;				//Driven by core logic
output 	PLLOUTCORE;				//PLL output to core logic
output	PLLOUTGLOBAL;	   			//PLL output to global network
input	EXTFEEDBACK;  				//Driven by core logic
input	[7:0] DYNAMICDELAY;  			//Driven by core logic
output	LOCK;					//Output of PLL
input	BYPASS;					//Driven by core logic
input	RESETB;					//Driven by core logic
input	LATCHINPUTVALUE; 			//iCEGate signal

//Test/Dynamic PLL configuration Pins
output	SDO;					//Output of PLL to core logic. 
input	SDI;					//Driven by core logic
input	SCLK;					//Driven by core logic

wire SPLLOUT1net;
wire SPLLOUT2net;

// Parameters 
parameter FEEDBACK_PATH = "SIMPLE";			//String  (simple, delay, phase_and_delay, external) 
parameter DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED"; 
parameter DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED"; 
parameter SHIFTREG_DIV_MODE = 2'b00; 			//0-->Divide by 4, 1-->Divide by 7, 3 -->Divide by 5
parameter FDA_FEEDBACK = 4'b0000; 			//Integer. 
parameter FDA_RELATIVE = 4'b0000; 			//Integer. 
parameter PLLOUT_SELECT = "GENCLK"; 			// 

//Use the Spreadsheet to populate the values below.
parameter DIVR = 4'b0000; 				//determine a good default value
parameter DIVF = 7'b0000000; 				//determine a good default value
parameter DIVQ = 3'b000; 				//determine a good default value
parameter FILTER_RANGE = 3'b000; 			//determine a good default value

parameter ENABLE_ICEGATE = 1'b0; 			//Additional cbits	
parameter TEST_MODE = 1'b0;				//TestMode parameter. Used for test/Dynamic PLL configuration.  
parameter EXTERNAL_DIVIDE_FACTOR = 1; 			//Not used by model. Added for PLL Config GUI.

generate

if(TEST_MODE==1) begin

	Sbt_DS_PLL40 instSbtSPLL (
		.CORE_REF_CLK (REFERENCECLK),
        	.PACKAGEPIN (),
		.EXTFEEDBACK (EXTFEEDBACK),  	
		.DYNAMICDELAY (DYNAMICDELAY),		
		.BYPASS (BYPASS),
		.RESETB (~RESETB),	
		.PLL_SCK(SCLK),
	        .PLL_SDI(SDI),
        	.PLL_SDO(SDO),
		.PLLOUT1 (SPLLOUT1net),	
		.PLLOUT2 (SPLLOUT2net),		
		.LOCK (LOCK)   	
	);	

	defparam instSbtSPLL.DIVR = DIVR;	
	defparam instSbtSPLL.DIVF = DIVF;
	defparam instSbtSPLL.DIVQ = DIVQ;
	defparam instSbtSPLL.FILTER_RANGE = FILTER_RANGE;
	defparam instSbtSPLL.FEEDBACK_PATH = FEEDBACK_PATH;
	defparam instSbtSPLL.DELAY_ADJUSTMENT_MODE_RELATIVE = DELAY_ADJUSTMENT_MODE_RELATIVE;
	defparam instSbtSPLL.DELAY_ADJUSTMENT_MODE_FEEDBACK = DELAY_ADJUSTMENT_MODE_FEEDBACK;
	defparam instSbtSPLL.SHIFTREG_DIV_MODE = SHIFTREG_DIV_MODE;
	defparam instSbtSPLL.FDA_RELATIVE = FDA_RELATIVE; 
	defparam instSbtSPLL.FDA_FEEDBACK = FDA_FEEDBACK; 
	defparam instSbtSPLL.PLLOUT_SELECT_PORTA = PLLOUT_SELECT;
	defparam instSbtSPLL.PLLOUT_SELECT_PORTB = "GENCLK";
	defparam instSbtSPLL.TEST_MODE = TEST_MODE;

end else begin

	SbtSPLL40 instSbtSPLL (
		.REFERENCECLK (REFERENCECLK),
		.EXTFEEDBACK (EXTFEEDBACK),  	
		.DYNAMICDELAY (DYNAMICDELAY),		
		.BYPASS (BYPASS),
		.RESETB (~RESETB),			
		.PLLOUT1 (SPLLOUT1net),	
		.PLLOUT2 (SPLLOUT2net),		
		.LOCK (LOCK)   	
	); 

	defparam instSbtSPLL.DIVR = DIVR;	
	defparam instSbtSPLL.DIVF = DIVF;
	defparam instSbtSPLL.DIVQ = DIVQ;
	defparam instSbtSPLL.FILTER_RANGE = FILTER_RANGE;
	defparam instSbtSPLL.FEEDBACK_PATH = FEEDBACK_PATH;
	defparam instSbtSPLL.DELAY_ADJUSTMENT_MODE_RELATIVE = DELAY_ADJUSTMENT_MODE_RELATIVE;
	defparam instSbtSPLL.DELAY_ADJUSTMENT_MODE_FEEDBACK = DELAY_ADJUSTMENT_MODE_FEEDBACK;
	defparam instSbtSPLL.SHIFTREG_DIV_MODE = SHIFTREG_DIV_MODE;
	defparam instSbtSPLL.FDA_RELATIVE = FDA_RELATIVE; 
	defparam instSbtSPLL.FDA_FEEDBACK = FDA_FEEDBACK; 
	defparam instSbtSPLL.PLLOUT_SELECT_PORTA = PLLOUT_SELECT;
	defparam instSbtSPLL.PLLOUT_SELECT_PORTB = "GENCLK";
	//defparam instSbtSPLL.TEST_MODE = TEST_MODE;
end	 
endgenerate			

assign PLLOUTCORE = ((ENABLE_ICEGATE != 0) && LATCHINPUTVALUE) ? PLLOUTCORE : SPLLOUT1net;
assign PLLOUTGLOBAL = ((ENABLE_ICEGATE != 0) && LATCHINPUTVALUE)  ? PLLOUTGLOBAL : SPLLOUT1net;

`ifdef TIMINGCHECK
specify
   (REFERENCECLK *> PLLOUTGLOBAL) = (1.0, 1.0);
   (REFERENCECLK *> PLLOUTCORE) = (1.0, 1.0);
   (SCLK *> SDO) = (1.0, 1.0);
   $setup(posedge SDI, posedge SCLK, 1.0);
   $setup(negedge SDI, posedge SCLK, 1.0);
   $setup(posedge SDI, negedge SCLK, 1.0);
   $setup(negedge SDI, negedge SCLK, 1.0);
   $hold(posedge SCLK, posedge SDI, 1.0);
   $hold(posedge SCLK, negedge SDI, 1.0);
   $hold(negedge SCLK, posedge SDI, 1.0);
   $hold(negedge SCLK, negedge SDI, 1.0);
endspecify
`endif
endmodule // SB_PLL40_CORE


////-----------------------------------------------------
//// ------------ SB_PLL40_PAD  -------------------------
////-----------------------------------------------------



`timescale 1ps/1ps
module SB_PLL40_PAD (
		PACKAGEPIN,		
		PLLOUTCORE,			//PLL output to core logic
		PLLOUTGLOBAL,	   		//PLL output to global network
		EXTFEEDBACK,  			//Driven by core logic
		DYNAMICDELAY,			//Driven by core logic
		LOCK,				//Output of PLL
		BYPASS,				//Driven by core logic
		RESETB,				//Driven by core logic
		SDI,				//Driven by core logic. Test Pin
		SDO,				//Output to RB Logic Tile. Test Pin
		SCLK,				//Driven by core logic. Test Pin
		LATCHINPUTVALUE 		//iCEGate signal
);
inout 	PACKAGEPIN;		
output 	PLLOUTCORE;				//PLL output to core logic
output	PLLOUTGLOBAL;	   			//PLL output to global network
input	EXTFEEDBACK;  				//Driven by core logic
input	[7:0] DYNAMICDELAY;  			//Driven by core logic
output	LOCK;					//Output of PLL
input	BYPASS;					//Driven by core logic
input	RESETB;					//Driven by core logic
input	LATCHINPUTVALUE; 			//iCEGate signal
//Test/Dynamic PLL configuration Pins
output	SDO;					//Output of PLL to core logic 
input	SDI;					//Driven by core logic
input	SCLK;					//Driven by core logic
wire SPLLOUT1net;

// Parameters 
parameter FEEDBACK_PATH = "SIMPLE";		//String  (simple, delay, phase_and_delay, external) 
parameter DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED"; 
parameter DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED"; 
parameter SHIFTREG_DIV_MODE = 2'b00; 		//0-->Divide by 4, 1-->Divide by 7, 3 -->Divide by 5
parameter FDA_FEEDBACK = 4'b0000; 		//Integer. 

parameter FDA_RELATIVE = 4'b0000; 		//Integer. 
parameter PLLOUT_SELECT = "GENCLK"; 		

//Use the Spreadsheet to populate the values below.
parameter DIVR = 4'b0000; 			//determine a good default value
parameter DIVF = 7'b0000000; 			//determine a good default value
parameter DIVQ = 3'b000; 			//determine a good default value
parameter FILTER_RANGE = 3'b000; 		//determine a good default value


parameter ENABLE_ICEGATE = 1'b0;		//Additional cbits
parameter TEST_MODE = 1'b0;			//Test Mode parameter.Used for test/Dynamic PLL configuration.  
parameter EXTERNAL_DIVIDE_FACTOR = 1; 		//Not used by model. Added for PLL Config GUI.	 


generate
if (TEST_MODE==1'b1) begin

	Sbt_DS_PLL40 instSbtSPLL (
		.CORE_REF_CLK (),
        	.PACKAGEPIN (PACKAGEPIN),
		.EXTFEEDBACK (EXTFEEDBACK),  	
		.DYNAMICDELAY (DYNAMICDELAY),		
		.BYPASS (BYPASS),
		.RESETB (~RESETB),	
		.PLL_SCK(SCLK),
	        .PLL_SDI(SDI),
        	.PLL_SDO(SDO),
		.PLLOUT1 (SPLLOUT1net),	
		.PLLOUT2 (SPLLOUT2net),		
		.LOCK (LOCK)   	

	);	   
	defparam instSbtSPLL.DIVR = DIVR;	
	defparam instSbtSPLL.DIVF = DIVF;
	defparam instSbtSPLL.DIVQ = DIVQ;
	defparam instSbtSPLL.FILTER_RANGE = FILTER_RANGE;
	defparam instSbtSPLL.FEEDBACK_PATH = FEEDBACK_PATH;
	defparam instSbtSPLL.DELAY_ADJUSTMENT_MODE_RELATIVE = DELAY_ADJUSTMENT_MODE_RELATIVE;
	defparam instSbtSPLL.DELAY_ADJUSTMENT_MODE_FEEDBACK = DELAY_ADJUSTMENT_MODE_FEEDBACK;
	defparam instSbtSPLL.SHIFTREG_DIV_MODE = SHIFTREG_DIV_MODE;
	defparam instSbtSPLL.FDA_RELATIVE = FDA_RELATIVE; 
	defparam instSbtSPLL.FDA_FEEDBACK = FDA_FEEDBACK; 
	defparam instSbtSPLL.PLLOUT_SELECT_PORTA = PLLOUT_SELECT;
	defparam instSbtSPLL.PLLOUT_SELECT_PORTB = "GENCLK";
	defparam instSbtSPLL.TEST_MODE = TEST_MODE;

end else begin

	SbtSPLL40 instSbtSPLL (
		.REFERENCECLK (PACKAGEPIN),
		.EXTFEEDBACK (EXTFEEDBACK),  	
		.DYNAMICDELAY (DYNAMICDELAY),		
		.BYPASS (BYPASS),
		.RESETB (~RESETB),			
		.PLLOUT1 (SPLLOUT1net),	
		.PLLOUT2 (SPLLOUT2net),		
		.LOCK (LOCK)   	
	);	  

	defparam instSbtSPLL.DIVR = DIVR;	
	defparam instSbtSPLL.DIVF = DIVF;
	defparam instSbtSPLL.DIVQ = DIVQ;
	defparam instSbtSPLL.FILTER_RANGE = FILTER_RANGE;
	defparam instSbtSPLL.FEEDBACK_PATH = FEEDBACK_PATH;
	defparam instSbtSPLL.DELAY_ADJUSTMENT_MODE_RELATIVE = DELAY_ADJUSTMENT_MODE_RELATIVE;
	defparam instSbtSPLL.DELAY_ADJUSTMENT_MODE_FEEDBACK = DELAY_ADJUSTMENT_MODE_FEEDBACK;
	defparam instSbtSPLL.SHIFTREG_DIV_MODE = SHIFTREG_DIV_MODE;
	defparam instSbtSPLL.FDA_RELATIVE = FDA_RELATIVE; 
	defparam instSbtSPLL.FDA_FEEDBACK = FDA_FEEDBACK; 
	defparam instSbtSPLL.PLLOUT_SELECT_PORTA = PLLOUT_SELECT;
	defparam instSbtSPLL.PLLOUT_SELECT_PORTB = "GENCLK";
	//defparam instSbtSPLL.TEST_MODE = TEST_MODE;

end

endgenerate

assign PLLOUTCORE = ((ENABLE_ICEGATE != 0) && LATCHINPUTVALUE) ? PLLOUTCORE : SPLLOUT1net;
assign PLLOUTGLOBAL = ((ENABLE_ICEGATE != 0) && LATCHINPUTVALUE)  ? PLLOUTGLOBAL : SPLLOUT1net;

`ifdef TIMINGCHECK
specify
   (PACKAGEPIN *> PLLOUTGLOBAL) = (1.0, 1.0);
   (PACKAGEPIN *> PLLOUTCORE) = (1.0, 1.0);
   (SCLK *> SDO) = (1.0, 1.0);
   $setup(posedge SDI, posedge SCLK, 1.0);
   $setup(negedge SDI, posedge SCLK, 1.0);
   $setup(posedge SDI, negedge SCLK, 1.0);
   $setup(negedge SDI, negedge SCLK, 1.0);
   $hold(posedge SCLK, posedge SDI, 1.0);
   $hold(posedge SCLK, negedge SDI, 1.0);
   $hold(negedge SCLK, posedge SDI, 1.0);
   $hold(negedge SCLK, negedge SDI, 1.0);
endspecify
`endif

endmodule // SB_PLL40_PAD

////-----------------------------------------------------
//// ------------ SB_PLL40_2_PAD  -----------------------
////-----------------------------------------------------

`timescale 1ps/1ps
module SB_PLL40_2_PAD (
		PACKAGEPIN,		
		PLLOUTCOREA,			//DIN0 output to core logic
		PLLOUTGLOBALA,	   		//GLOBALOUTPUTBUFFER
	        PLLOUTCOREB,			//PLL output to core logic
		PLLOUTGLOBALB,	   		//PLL output to global network
		EXTFEEDBACK,  			//Driven by core logic
		DYNAMICDELAY,			//Driven by core logic
		LOCK,				//Output of PLL
		BYPASS,				//Driven by core logic
		RESETB,				//Driven by core logic
		SDI,				//Driven by core logic. Test Pin
		SDO,				//Output to RB Logic Tile. Test Pin
		SCLK,				//Driven by core logic. Test Pin
		LATCHINPUTVALUE 		//iCEGate signal
);
inout 	PACKAGEPIN;		
output  PLLOUTCOREA;				//PLL output to core logic
output	PLLOUTGLOBALA;	   			//PLL output to global network
output  PLLOUTCOREB;				//PLL output to core logic
output	PLLOUTGLOBALB;	   			//PLL output to global network
input	EXTFEEDBACK;  				//Driven by core logic
input	[7:0] DYNAMICDELAY;  			//Driven by core logic
output	LOCK;					//Output of PLL
input	BYPASS;					//Driven by core logic
input	RESETB;					//Driven by core logic
input	LATCHINPUTVALUE; 			//iCEGate signal
//Test/Dynamic PLL configuration Pins
output	SDO;					//Output of PLL to core logic. 
input	SDI;					//Driven by core logic
input	SCLK;					//Driven by core logic
wire SPLLOUT2net;

// Parameters 
parameter FEEDBACK_PATH = "SIMPLE";			//String  (simple, delay, phase_and_delay, external) 
parameter DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED"; 
parameter DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED"; 
parameter SHIFTREG_DIV_MODE = 2'b00; 			//0-->Divide by 4, 1-->Divide by 7, 3 -->Divide by 5
parameter FDA_FEEDBACK = 4'b0000; 			//Integer. 

//Output 
parameter FDA_RELATIVE = 4'b0000; 			//Integer. 
parameter PLLOUT_SELECT_PORTB = "GENCLK"; 		

//Use the Spreadsheet to populate the values below.
parameter DIVR = 4'b0000; 				//determine a good default value
parameter DIVF = 7'b0000000; 				//determine a good default value
parameter DIVQ = 3'b000; 				//determine a good default value
parameter FILTER_RANGE = 3'b000; 			//determine a good default value


parameter ENABLE_ICEGATE_PORTA = 1'b0;			//Additional cbits
parameter ENABLE_ICEGATE_PORTB = 1'b0;
parameter TEST_MODE = 1'b0;				//Test Mode parameter.Used for test/Dynamic PLL configuration.  
parameter EXTERNAL_DIVIDE_FACTOR = 1; 			//Not used by model. Added for PLL Config GUI.

generate

if(TEST_MODE==1'b1) begin

	Sbt_DS_PLL40 instSbtSPLL (
		.CORE_REF_CLK (),
        	.PACKAGEPIN (PACKAGEPIN),
		.EXTFEEDBACK (EXTFEEDBACK),  	
		.DYNAMICDELAY (DYNAMICDELAY),		
		.BYPASS (BYPASS),
		.RESETB (~RESETB),	
		.PLL_SCK(SCLK),
	        .PLL_SDI(SDI),
        	.PLL_SDO(SDO),
		.PLLOUT1 (SPLLOUT1net),	
		.PLLOUT2 (SPLLOUT2net),		
		.LOCK (LOCK)   	

	);	 
	defparam instSbtSPLL.DIVR = DIVR;	
	defparam instSbtSPLL.DIVF = DIVF;
	defparam instSbtSPLL.DIVQ = DIVQ;
	defparam instSbtSPLL.FILTER_RANGE = FILTER_RANGE;
	defparam instSbtSPLL.FEEDBACK_PATH = FEEDBACK_PATH;
	defparam instSbtSPLL.DELAY_ADJUSTMENT_MODE_RELATIVE = DELAY_ADJUSTMENT_MODE_RELATIVE;
	defparam instSbtSPLL.DELAY_ADJUSTMENT_MODE_FEEDBACK = DELAY_ADJUSTMENT_MODE_FEEDBACK;
	defparam instSbtSPLL.SHIFTREG_DIV_MODE = SHIFTREG_DIV_MODE;
	defparam instSbtSPLL.FDA_RELATIVE = FDA_RELATIVE; 
	defparam instSbtSPLL.FDA_FEEDBACK = FDA_FEEDBACK; 
	defparam instSbtSPLL.PLLOUT_SELECT_PORTA = "GENCLK";
	defparam instSbtSPLL.PLLOUT_SELECT_PORTB = PLLOUT_SELECT_PORTB;
	defparam instSbtSPLL.TEST_MODE = TEST_MODE;

end  else begin

	SbtSPLL40 instSbtSPLL (
		.REFERENCECLK (PACKAGEPIN),
		.EXTFEEDBACK (EXTFEEDBACK),  	
		.DYNAMICDELAY (DYNAMICDELAY),		
		.BYPASS (BYPASS),
		.RESETB (~RESETB),			
		.PLLOUT1 (SPLLOUT1net),	
		.PLLOUT2 (SPLLOUT2net),		
		.LOCK (LOCK)   	
	);	
	defparam instSbtSPLL.DIVR = DIVR;	
	defparam instSbtSPLL.DIVF = DIVF;
	defparam instSbtSPLL.DIVQ = DIVQ;
	defparam instSbtSPLL.FILTER_RANGE = FILTER_RANGE;
	defparam instSbtSPLL.FEEDBACK_PATH = FEEDBACK_PATH;
	defparam instSbtSPLL.DELAY_ADJUSTMENT_MODE_RELATIVE = DELAY_ADJUSTMENT_MODE_RELATIVE;
	defparam instSbtSPLL.DELAY_ADJUSTMENT_MODE_FEEDBACK = DELAY_ADJUSTMENT_MODE_FEEDBACK;
	defparam instSbtSPLL.SHIFTREG_DIV_MODE = SHIFTREG_DIV_MODE;
	defparam instSbtSPLL.FDA_RELATIVE = FDA_RELATIVE; 
	defparam instSbtSPLL.FDA_FEEDBACK = FDA_FEEDBACK; 
	defparam instSbtSPLL.PLLOUT_SELECT_PORTA = "GENCLK";
	defparam instSbtSPLL.PLLOUT_SELECT_PORTB = PLLOUT_SELECT_PORTB;
	//defparam instSbtSPLL.TEST_MODE = TEST_MODE;
end

endgenerate

assign PLLOUTCOREA = ((ENABLE_ICEGATE_PORTA != 0) && LATCHINPUTVALUE) ? PLLOUTCOREA : PACKAGEPIN;
assign PLLOUTGLOBALA = ((ENABLE_ICEGATE_PORTA != 0) && LATCHINPUTVALUE)  ? PLLOUTGLOBALA : PACKAGEPIN;
assign PLLOUTCOREB = ((ENABLE_ICEGATE_PORTB != 0) && LATCHINPUTVALUE) ? PLLOUTCOREB : SPLLOUT2net;
assign PLLOUTGLOBALB = ((ENABLE_ICEGATE_PORTB != 0) && LATCHINPUTVALUE)  ? PLLOUTGLOBALB : SPLLOUT2net;

`ifdef TIMINGCHECK
specify
   (PACKAGEPIN *> PLLOUTGLOBALA) = (1.0, 1.0);
   (PACKAGEPIN *> PLLOUTCOREA) = (1.0, 1.0);
   (PACKAGEPIN *> PLLOUTGLOBALB) = (1.0, 1.0);
   (PACKAGEPIN *> PLLOUTCOREB) = (1.0, 1.0);
   (SCLK *> SDO) = (1.0, 1.0);
   $setup(posedge SDI, posedge SCLK, 1.0);
   $setup(negedge SDI, posedge SCLK, 1.0);
   $setup(posedge SDI, negedge SCLK, 1.0);
   $setup(negedge SDI, negedge SCLK, 1.0);
   $hold(posedge SCLK, posedge SDI, 1.0);
   $hold(posedge SCLK, negedge SDI, 1.0);
   $hold(negedge SCLK, posedge SDI, 1.0);
   $hold(negedge SCLK, negedge SDI, 1.0);

endspecify
`endif

endmodule // SB_PLL40_2_PAD

////-----------------------------------------------------
//// ------------ SB_PLL40_2F_CORE ----------------------
////-----------------------------------------------------

`timescale 1ps/1ps
module SB_PLL40_2F_CORE (
		REFERENCECLK,			//Driven by core logic
		PLLOUTCOREA,			//DIN0 output to core logic
		PLLOUTGLOBALA,	   		//GLOBALOUTPUTBUFFER
	        PLLOUTCOREB,			//PLL output to core logic
		PLLOUTGLOBALB,	   		//PLL output to global network
		EXTFEEDBACK,  			//Driven by core logic
		DYNAMICDELAY,			//Driven by core logic
		LOCK,				//Output of PLL
		BYPASS,				//Driven by core logic
		RESETB,				//Driven by core logic
		SDI,				//Driven by core logic. Test Pin
		SDO,				//Output to RB Logic Tile. Test Pin
		SCLK,				//Driven by core logic. Test Pin
		LATCHINPUTVALUE 		//iCEGate signal
);
input 	REFERENCECLK;				//Driven by core logic
output  PLLOUTCOREA;				//PLL output to core logic
output	PLLOUTGLOBALA;	   			//PLL output to global network
output  PLLOUTCOREB;				//PLL output to core logic
output	PLLOUTGLOBALB;	   			//PLL output to global network
input	EXTFEEDBACK;  				//Driven by core logic
input	[7:0] DYNAMICDELAY;  			//Driven by core logic
output	LOCK;					//Output of PLL
input	BYPASS;					//Driven by core logic
input	RESETB;					//Driven by core logic
input	LATCHINPUTVALUE; 			//iCEGate signal
//Test/Dynamic PLL configuration Pins
output	SDO;					//Output of PLL
input	SDI;					//Driven by core logic
input	SCLK;					//Driven by core logic

wire SPLLOUT1net;
wire SPLLOUT2net;

// Parameters 
parameter FEEDBACK_PATH = "SIMPLE";			//String  (simple, delay, phase_and_delay, external) 
parameter DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED"; 
parameter DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED"; 
parameter SHIFTREG_DIV_MODE = 2'b00; 			//0-->Divide by 4, 1-->Divide by 7, 3 -->Divide by 5
parameter FDA_FEEDBACK = 4'b0000; 			//Integer. 
parameter FDA_RELATIVE = 4'b0000; 			//Integer. 
parameter PLLOUT_SELECT_PORTA = "GENCLK"; 		//
parameter PLLOUT_SELECT_PORTB = "GENCLK"; 		//
//Use the Spreadsheet to populate the values below.
parameter DIVR = 4'b0000; 				//determine a good default value
parameter DIVF = 7'b0000000; 				//determine a good default value
parameter DIVQ = 3'b000; 				//determine a good default value
parameter FILTER_RANGE = 3'b000; 			//determine a good default value						
parameter ENABLE_ICEGATE_PORTA = 1'b0;			//Additional cbits
parameter ENABLE_ICEGATE_PORTB = 1'b0;
parameter TEST_MODE = 1'b0;				//Test Mode parameter.Used for test/Dynamic PLL configuration.
parameter EXTERNAL_DIVIDE_FACTOR = 1; 			//Not used by model. Added for PLL Config GUI.
generate
if(TEST_MODE==1) begin

	Sbt_DS_PLL40 instSbtSPLL (
		.CORE_REF_CLK (REFERENCECLK),
	        .PACKAGEPIN (),
		.EXTFEEDBACK (EXTFEEDBACK),  	
		.DYNAMICDELAY (DYNAMICDELAY),		
		.BYPASS (BYPASS),
		.RESETB (~RESETB),	
		.PLL_SCK(SCLK),
        	.PLL_SDI(SDI),
        	.PLL_SDO(SDO),
		.PLLOUT1 (SPLLOUT1net),	
		.PLLOUT2 (SPLLOUT2net),		
		.LOCK (LOCK)   	
	);	
	defparam instSbtSPLL.DIVR = DIVR;	
	defparam instSbtSPLL.DIVF = DIVF;
	defparam instSbtSPLL.DIVQ = DIVQ;
	defparam instSbtSPLL.FILTER_RANGE = FILTER_RANGE;
	defparam instSbtSPLL.FEEDBACK_PATH = FEEDBACK_PATH;
	defparam instSbtSPLL.DELAY_ADJUSTMENT_MODE_RELATIVE = DELAY_ADJUSTMENT_MODE_RELATIVE;
	defparam instSbtSPLL.DELAY_ADJUSTMENT_MODE_FEEDBACK = DELAY_ADJUSTMENT_MODE_FEEDBACK;
	defparam instSbtSPLL.SHIFTREG_DIV_MODE = SHIFTREG_DIV_MODE;
	defparam instSbtSPLL.FDA_RELATIVE = FDA_RELATIVE; 
	defparam instSbtSPLL.FDA_FEEDBACK = FDA_FEEDBACK; 
	defparam instSbtSPLL.PLLOUT_SELECT_PORTA = PLLOUT_SELECT_PORTA;
	defparam instSbtSPLL.PLLOUT_SELECT_PORTB = PLLOUT_SELECT_PORTB;
	defparam instSbtSPLL.TEST_MODE = TEST_MODE;

end else begin
	SbtSPLL40 instSbtSPLL (
		.REFERENCECLK (REFERENCECLK),
		.EXTFEEDBACK (EXTFEEDBACK),  	
		.DYNAMICDELAY (DYNAMICDELAY),		
		.BYPASS (BYPASS),
		.RESETB (~RESETB),			
		.PLLOUT1 (SPLLOUT1net),	
		.PLLOUT2 (SPLLOUT2net),		
		.LOCK (LOCK)   	

	);
	defparam instSbtSPLL.DIVR = DIVR;	
	defparam instSbtSPLL.DIVF = DIVF;
	defparam instSbtSPLL.DIVQ = DIVQ;
	defparam instSbtSPLL.FILTER_RANGE = FILTER_RANGE;
	defparam instSbtSPLL.FEEDBACK_PATH = FEEDBACK_PATH;
	defparam instSbtSPLL.DELAY_ADJUSTMENT_MODE_RELATIVE = DELAY_ADJUSTMENT_MODE_RELATIVE;
	defparam instSbtSPLL.DELAY_ADJUSTMENT_MODE_FEEDBACK = DELAY_ADJUSTMENT_MODE_FEEDBACK;
	defparam instSbtSPLL.SHIFTREG_DIV_MODE = SHIFTREG_DIV_MODE;
	defparam instSbtSPLL.FDA_RELATIVE = FDA_RELATIVE; 
	defparam instSbtSPLL.FDA_FEEDBACK = FDA_FEEDBACK; 
	defparam instSbtSPLL.PLLOUT_SELECT_PORTA = PLLOUT_SELECT_PORTA;
	defparam instSbtSPLL.PLLOUT_SELECT_PORTB = PLLOUT_SELECT_PORTB;

end	 
endgenerate	

assign PLLOUTCOREA = ((ENABLE_ICEGATE_PORTA != 0) && LATCHINPUTVALUE) ? PLLOUTCOREA : SPLLOUT1net;
assign PLLOUTGLOBALA = ((ENABLE_ICEGATE_PORTA != 0) && LATCHINPUTVALUE)  ? PLLOUTGLOBALA : SPLLOUT1net;
assign PLLOUTCOREB = ((ENABLE_ICEGATE_PORTB != 0) && LATCHINPUTVALUE) ? PLLOUTCOREB : SPLLOUT2net;
assign PLLOUTGLOBALB = ((ENABLE_ICEGATE_PORTB != 0) && LATCHINPUTVALUE)  ? PLLOUTGLOBALB : SPLLOUT2net;

`ifdef TIMINGCHECK
specify
   (REFERENCECLK *> PLLOUTGLOBALA) = (1.0, 1.0);
   (REFERENCECLK *> PLLOUTCOREA) = (1.0, 1.0);
   (REFERENCECLK *> PLLOUTGLOBALB) = (1.0, 1.0);
   (REFERENCECLK *> PLLOUTCOREB) = (1.0, 1.0);
   (SCLK *> SDO) = (1.0, 1.0);
   $setup(posedge SDI, posedge SCLK, 1.0);
   $setup(negedge SDI, posedge SCLK, 1.0);
   $setup(posedge SDI, negedge SCLK, 1.0);
   $setup(negedge SDI, negedge SCLK, 1.0);
   $hold(posedge SCLK, posedge SDI, 1.0);
   $hold(posedge SCLK, negedge SDI, 1.0);
   $hold(negedge SCLK, posedge SDI, 1.0);
   $hold(negedge SCLK, negedge SDI, 1.0);
endspecify
`endif

endmodule // SB_PLL40_2F_CORE

////-----------------------------------------------------
//// ------------ SB_PLL40_2F_PAD  ----------------------
////-----------------------------------------------------


`timescale 1ps/1ps
module SB_PLL40_2F_PAD (
		PACKAGEPIN,		
		PLLOUTCOREA,			//DIN0 output to core logic
		PLLOUTGLOBALA,	   		//PLL output to global network
        	PLLOUTCOREB,			//PLL output to core logic
		PLLOUTGLOBALB,	   		//PLL output to global network
		EXTFEEDBACK,  			//Driven by core logic
		DYNAMICDELAY,			//Driven by core logic
		LOCK,				//Output of PLL
		BYPASS,				//Driven by core logic
		RESETB,				//Driven by core logic
		SDI,				//Driven by core logic. Test Pin
		SDO,				//Output to RB Logic Tile. Test Pin
		SCLK,				//Driven by core logic. Test Pin
		LATCHINPUTVALUE 		//iCEGate signal
);

inout 	PACKAGEPIN;		
output  PLLOUTCOREA;				//PLL output to core logic
output	PLLOUTGLOBALA;	   			//PLL output to global network
output  PLLOUTCOREB;				//PLL output to core logic
output	PLLOUTGLOBALB;	   			//PLL output to global network
input	EXTFEEDBACK;  				//Driven by core logic
input	[7:0] DYNAMICDELAY;  			//Driven by core logic
output	LOCK;					//Output of PLL
input	BYPASS;					//Driven by core logic
input	RESETB;					//Driven by core logic
input	LATCHINPUTVALUE; 			//iCEGate signal
//Test/Dynamic PLL configuration Pins 
output	SDO;					//Output of PLL
input	SDI;					//Driven by core logic
input	SCLK;					//Driven by core logic
wire SPLLOUT1net;
wire SPLLOUT2net;

// Parameters 
parameter FEEDBACK_PATH = "SIMPLE";		//String  (simple, delay, phase_and_delay, external) 
parameter DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED"; 
parameter DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED"; 
parameter SHIFTREG_DIV_MODE = 2'b00; 		//0-->Divide by 4, 1-->Divide by 7, 3 -->Divide by 5
parameter FDA_FEEDBACK = 4'b0000; 		//Integer. 
parameter FDA_RELATIVE = 4'b0000; 		//Integer. 
parameter PLLOUT_SELECT_PORTA = "GENCLK"; 	//
parameter PLLOUT_SELECT_PORTB = "GENCLK"; 	//
//Use the Spreadsheet to populate the values below.
parameter DIVR = 4'b0000; 			//determine a good default value
parameter DIVF = 7'b0000000; 			//determine a good default value
parameter DIVQ = 3'b000; 			//determine a good default value
parameter FILTER_RANGE = 3'b000; 		//determine a good default value
parameter ENABLE_ICEGATE_PORTA = 1'b0;		//Additional cbits
parameter ENABLE_ICEGATE_PORTB = 1'b0;
parameter TEST_MODE = 1'b0;			//Test Mode parameter.Used for test/Dynamic PLL configuration.
parameter EXTERNAL_DIVIDE_FACTOR = 1; 		//Not used by model. Added for PLL Config GUI.

generate
if(TEST_MODE==1) begin
	Sbt_DS_PLL40 instSbtSPLL (
		.CORE_REF_CLK (),
	        .PACKAGEPIN (PACKAGEPIN),
		.EXTFEEDBACK (EXTFEEDBACK),  	
		.DYNAMICDELAY (DYNAMICDELAY),		
		.BYPASS (BYPASS),
		.RESETB (~RESETB),	
		.PLL_SCK(SCLK),
        	.PLL_SDI(SDI),
        	.PLL_SDO(SDO),
		.PLLOUT1 (SPLLOUT1net),	
		.PLLOUT2 (SPLLOUT2net),		
		.LOCK (LOCK)   
		);	

	defparam instSbtSPLL.DIVR = DIVR;	
	defparam instSbtSPLL.DIVF = DIVF;
	defparam instSbtSPLL.DIVQ = DIVQ;
	defparam instSbtSPLL.FILTER_RANGE = FILTER_RANGE;
	defparam instSbtSPLL.FEEDBACK_PATH = FEEDBACK_PATH;
	defparam instSbtSPLL.DELAY_ADJUSTMENT_MODE_RELATIVE = DELAY_ADJUSTMENT_MODE_RELATIVE;
	defparam instSbtSPLL.DELAY_ADJUSTMENT_MODE_FEEDBACK = DELAY_ADJUSTMENT_MODE_FEEDBACK;
	defparam instSbtSPLL.SHIFTREG_DIV_MODE = SHIFTREG_DIV_MODE;
	defparam instSbtSPLL.FDA_RELATIVE = FDA_RELATIVE; 
	defparam instSbtSPLL.FDA_FEEDBACK = FDA_FEEDBACK; 
	defparam instSbtSPLL.PLLOUT_SELECT_PORTA = PLLOUT_SELECT_PORTA;
	defparam instSbtSPLL.PLLOUT_SELECT_PORTB = PLLOUT_SELECT_PORTB;
	defparam instSbtSPLL.TEST_MODE = TEST_MODE;

end else begin
	SbtSPLL40 instSbtSPLL (
		.REFERENCECLK (PACKAGEPIN),
		.EXTFEEDBACK (EXTFEEDBACK),  	
		.DYNAMICDELAY (DYNAMICDELAY),		
		.BYPASS (BYPASS),
		.RESETB (~RESETB),			
		.PLLOUT1 (SPLLOUT1net),	
		.PLLOUT2 (SPLLOUT2net),		
		.LOCK (LOCK)   	
	);

	defparam instSbtSPLL.DIVR = DIVR;	
	defparam instSbtSPLL.DIVF = DIVF;
	defparam instSbtSPLL.DIVQ = DIVQ;
	defparam instSbtSPLL.FILTER_RANGE = FILTER_RANGE;
	defparam instSbtSPLL.FEEDBACK_PATH = FEEDBACK_PATH;
	defparam instSbtSPLL.DELAY_ADJUSTMENT_MODE_RELATIVE = DELAY_ADJUSTMENT_MODE_RELATIVE;
	defparam instSbtSPLL.DELAY_ADJUSTMENT_MODE_FEEDBACK = DELAY_ADJUSTMENT_MODE_FEEDBACK;
	defparam instSbtSPLL.SHIFTREG_DIV_MODE = SHIFTREG_DIV_MODE;
	defparam instSbtSPLL.FDA_RELATIVE = FDA_RELATIVE; 
	defparam instSbtSPLL.FDA_FEEDBACK = FDA_FEEDBACK; 
	defparam instSbtSPLL.PLLOUT_SELECT_PORTA = PLLOUT_SELECT_PORTA;
	defparam instSbtSPLL.PLLOUT_SELECT_PORTB = PLLOUT_SELECT_PORTB;

end	 
endgenerate	

assign PLLOUTCOREA = ((ENABLE_ICEGATE_PORTA != 0) && LATCHINPUTVALUE) ? PLLOUTCOREA : SPLLOUT1net;
assign PLLOUTGLOBALA = ((ENABLE_ICEGATE_PORTA != 0) && LATCHINPUTVALUE)  ? PLLOUTGLOBALA : SPLLOUT1net;
assign PLLOUTCOREB = ((ENABLE_ICEGATE_PORTB != 0) && LATCHINPUTVALUE) ? PLLOUTCOREB : SPLLOUT2net;
assign PLLOUTGLOBALB = ((ENABLE_ICEGATE_PORTB != 0) && LATCHINPUTVALUE)  ? PLLOUTGLOBALB : SPLLOUT2net;

 
`ifdef TIMINGCHECK
specify
   (PACKAGEPIN *> PLLOUTGLOBALA) = (1.0, 1.0);
   (PACKAGEPIN *> PLLOUTCOREA) = (1.0, 1.0);
   (PACKAGEPIN *> PLLOUTGLOBALB) = (1.0, 1.0);
   (PACKAGEPIN *> PLLOUTCOREB) = (1.0, 1.0);
   (SCLK *> SDO) = (1.0, 1.0);
   $setup(posedge SDI, posedge SCLK, 1.0);
   $setup(negedge SDI, posedge SCLK, 1.0);
   $setup(posedge SDI, negedge SCLK, 1.0);
   $setup(negedge SDI, negedge SCLK, 1.0);
   $hold(posedge SCLK, posedge SDI, 1.0);
   $hold(posedge SCLK, negedge SDI, 1.0);
   $hold(negedge SCLK, posedge SDI, 1.0);
   $hold(negedge SCLK, negedge SDI, 1.0);
endspecify
`endif

endmodule // SB_PLL40_2F_PAD

////-----------------------------------------------------
//// ------------ SB_MIPI_RX_2LANE ----------------------
////-----------------------------------------------------


`timescale 1ps/1ps
module    SB_MIPI_RX_2LANE(
  ENPDESER,
  PU,
  DP0,
  DN0,
  D0RXHSEN,
  D0DTXLPP,
  D0DTXLPN,
  D0TXLPEN,
  D0DRXLPP,
  D0DRXLPN,
  D0RXLPEN,
  D0DCDP,
  D0DCDN,
  D0CDEN,
  D0HSDESEREN,
  D0HSRXDATA,
  D0HSBYTECLKD,
  D0SYNC,
  D0ERRSYNC,
  D0NOSYNC,
  DP1,
  DN1,
  D1RXHSEN,
  D1DRXLPP,
  D1DRXLPN,
  D1RXLPEN,
  D1HSDESEREN,
  D1HSRXDATA,
  D1SYNC,
  D1ERRSYNC,
  D1NOSYNC,
  CKP,
  CKN,
  CLKRXHSEN,
  CLKDRXLPP,
  CLKDRXLPN,
  CLKRXLPEN,
  CLKHSBYTE
  );

// Device pins are DP1,DN1,DP0,DN0,CKP,CKN

//Common Interface Pins
input         ENPDESER;
input 			     PU;
//input				     LBEN;


// DATA0 Interface pins
input				     DP0;
input				     DN0;
input				     D0RXHSEN;
//input				     D0RXHSTHDB;
input 			     D0DTXLPP;
input 			     D0DTXLPN;
input  			    D0TXLPEN;
output 			    D0DRXLPP;
output  			   D0DRXLPN;
input 			     D0RXLPEN;
output 			    D0DCDP;
output			     D0DCDN;
input 			     D0CDEN;
input				     D0HSDESEREN;
output  [7:0]	D0HSRXDATA;
output 			    D0HSBYTECLKD;
output  			   D0SYNC;
output  			   D0ERRSYNC;
output 			    D0NOSYNC;
//output        D0DRXHS;

// DATA1 Interface Pins
input  			    DP1;
input  			    DN1;
input  			    D1RXHSEN;
//input  			    D1RXHSTHDB;
output  			   D1DRXLPP;
output  			   D1DRXLPN;
input  			    D1RXLPEN;
//output  			   D1DCDP;
//output  			   D1DCDN;
//input  			    D1CDEN;
input  			    D1HSDESEREN;
output  [7:0] D1HSRXDATA;
output  			   D1SYNC;
output  			   D1ERRSYNC;
output  			   D1NOSYNC;
//output        D1DRXHS;


// CLOCK Interface Pins
input  			    CKP;
input  			    CKN;
input  			    CLKRXHSEN;
//input  			    CLKRXHSTHDB;
output  			   CLKDRXLPP;
output  			   CLKDRXLPN;
input  			    CLKRXLPEN;
//output  			   CLKDCDP;
//output  			   CLKDCDN;
//input  			    CLKCDEN;

output        CLKHSBYTE;
//output        CLKDRXHS;

X105DSI_RX                  u_mipi_slave_analog(
// Power and Ground Pins
  .VDDA                   (1'b1),
  .VSSA                   (1'b0),
  .DVSS                   (1'b0),
 // Common Interface pins 
  .ENP_DESER              (ENPDESER),
  .PD                     (~PU),
 //Data0 Interface pins
  .DP0                    (DP0),
  .DN0                    (DN0),
  .D0_RXHSEN              (D0RXHSEN),
  .D0_DTXLPP              (D0DTXLPP),
  .D0_DTXLPN              (D0DTXLPN),
  .D0_TXLPEN              (D0TXLPEN),
  .D0_DRXLPP              (D0DRXLPP),
  .D0_DRXLPN              (D0DRXLPN),
  .D0_RXLPEN              (D0RXLPEN),
  .D0_DCDP                (D0DCDP),
  .D0_DCDN                (D0DCDN),
  .D0_CDEN                (D0CDEN),
  .D0_HS_DESER_EN         (D0HSDESEREN),
  .D0_HSRX_DATA           (D0HSRXDATA),
  .D0_HS_BYTE_CLKD        (D0HSBYTECLKD),
  .D0_SYNC                (D0SYNC),
  .D0_ERRSYNC             (D0ERRSYNC),
  .D0_NOSYNC              (D0NOSYNC),
 // DATA1 Interface pins
  .DP1                    (DP1),
  .DN1                    (DN1),
  .D1_RXHSEN              (D1RXHSEN),
  .D1_DRXLPP              (D1DRXLPP),
  .D1_DRXLPN              (D1DRXLPN),
  .D1_RXLPEN              (D1RXLPEN),
  .D1_HS_DESER_EN         (D1HSDESEREN),
  .D1_HSRX_DATA           (D1HSRXDATA),
  .D1_SYNC                (D1SYNC),
  .D1_ERRSYNC             (D1ERRSYNC),
  .D1_NOSYNC              (D1NOSYNC),
 // CLOCK Interface pins
  .CKP                    (CKP),
  .CKN                    (CKN),
  .CLK_RXHSEN             (CLKRXHSEN),
  .CLK_DRXLPP             (CLKDRXLPP),
  .CLK_DRXLPN             (CLKDRXLPN),
  .CLK_RXLPEN             (CLKRXLPEN),
  .CLK_HS_BYTE            (CLKHSBYTE)
  );

`ifdef TIMINGCHECK
specify
    //Data0 Lane tp & tCQ 
   (DP0 *> D0DRXLPP) = (1.0, 1.0);
   (DN0 *> D0DRXLPN) = (1.0, 1.0);	
   (DP0 *> D0DCDP  ) = (1.0, 1.0);	  
   (DN0 *> D0DCDN  ) = (1.0, 1.0); 
   (CKP *> D0HSRXDATA[0]) = (1.0, 1.0);	
   (CKP *> D0HSRXDATA[1]) = (1.0, 1.0);	
   (CKP *> D0HSRXDATA[2]) = (1.0, 1.0);	
   (CKP *> D0HSRXDATA[3]) = (1.0, 1.0);	
   (CKP *> D0HSRXDATA[4]) = (1.0, 1.0);	
   (CKP *> D0HSRXDATA[5]) = (1.0, 1.0);	
   (CKP *> D0HSRXDATA[6]) = (1.0, 1.0);	
   (CKP *> D0HSRXDATA[7]) = (1.0, 1.0);	
   (CKP *> D0HSBYTECLKD ) = (1.0, 1.0);	 
    //Data1 Lane tp & tCQ 
   (DP1 *> D1DRXLPP) = (1.0, 1.0);
   (DN1 *> D1DRXLPN) = (1.0, 1.0);	
   (CKP *> D1HSRXDATA[0]) = (1.0, 1.0);	
   (CKP *> D1HSRXDATA[1]) = (1.0, 1.0);	
   (CKP *> D1HSRXDATA[2]) = (1.0, 1.0);	
   (CKP *> D1HSRXDATA[3]) = (1.0, 1.0);	
   (CKP *> D1HSRXDATA[4]) = (1.0, 1.0);	
   (CKP *> D1HSRXDATA[5]) = (1.0, 1.0);	
   (CKP *> D1HSRXDATA[6]) = (1.0, 1.0);	
   (CKP *> D1HSRXDATA[7]) = (1.0, 1.0);	
   //Clk Lane tp & tCQ 			  
   (CKP  *> CLKDRXLPP ) = (1.0, 1.0);
   (CKN  *> CLKDRXLPN ) = (1.0, 1.0);
   (CKP  *> CLKHSBYTE) = (1.0, 1.0);
   // Data0 Lane setup-hold cheks 
   $setup(posedge DP0, posedge CKP, 1.0);
   $setup(negedge DP0, posedge CKP, 1.0);
   $hold (posedge CKP, posedge DP0, 1.0);
   $hold (posedge CKP, negedge DP0, 1.0);   
   $setup(posedge DP0, negedge CKP, 1.0);
   $setup(negedge DP0, negedge CKP, 1.0);
   $hold (negedge CKP, posedge DP0, 1.0);
   $hold (negedge CKP, negedge DP0, 1.0);
   
   $setup(posedge DN0, posedge CKP, 1.0);
   $setup(negedge DN0, posedge CKP, 1.0);
   $hold (posedge CKP, posedge DN0, 1.0);
   $hold (posedge CKP, negedge DN0, 1.0);   
   $setup(posedge DN0, negedge CKP, 1.0);
   $setup(negedge DN0, negedge CKP, 1.0);
   $hold (negedge CKP, posedge DN0, 1.0);
   $hold (negedge CKP, negedge DN0, 1.0);
   // Data 1 Lane setup-hold checks  
   $setup(posedge DP1, posedge CKP, 1.0);
   $setup(negedge DP1, posedge CKP, 1.0);
   $hold (posedge CKP, posedge DP1, 1.0);
   $hold (posedge CKP, negedge DP1, 1.0);   
   $setup(posedge DP1, negedge CKP, 1.0);
   $setup(negedge DP1, negedge CKP, 1.0);
   $hold (negedge CKP, posedge DP1, 1.0);
   $hold (negedge CKP, negedge DP1, 1.0);  
   
   $setup(posedge DN1, posedge CKP, 1.0);
   $setup(negedge DN1, posedge CKP, 1.0);
   $hold (posedge CKP, posedge DN1, 1.0);
   $hold (posedge CKP, negedge DN1, 1.0);   
   $setup(posedge DN1, negedge CKP, 1.0);
   $setup(negedge DN1, negedge CKP, 1.0);
   $hold (negedge CKP, posedge DN1, 1.0);
   $hold (negedge CKP, negedge DN1, 1.0);      
endspecify
`endif   
  
endmodule

`timescale 1ps/1ps
 
module SB_TMDS_deserializer(
                                //TMDS input interface
  input TMDSch0p,             //TMDS ch 0 differential input pos
  input TMDSch0n,             //TMDS ch 0 differential input neg
  input TMDSch1p,             //TMDS ch 1 differential input pos
  input TMDSch1n,             //TMDS ch 1 differential input neg
  input TMDSch2p,             //TMDS ch 2 differential input pos
  input TMDSch2n,             //TMDS ch 2 differential input neg
  input TMDSclkp,             //TMDS clock differential input pos
  input TMDSclkn,             //TMDS clock differential input neg
                                
                                //Receive controller interface
  input RSTNdeser,             //Reset deserailzier logics- active low
  input RSTNpll,               //Reset deserializer PLL- active low
  input EN,                     //Enable deserializer- active high
  input [3:0] PHASELch0,       //Clock phase delay compensation select for ch 0
  input [3:0] PHASELch1,       //Clock phase delay compensation select for ch 1
  input [3:0] PHASELch2,       //Clock phase delay compensation select for ch 2
  output PLLlock,              //PLL lock signal- active high
  output PLLOUTGLOBALclkx1,    //PLL output on global n/w 
  output PLLOUTCOREclkx1,    	//PLL output on global n/w 
  output PLLOUTGLOBALclkx5,    //PLL output on global n/w 
  output PLLOUTCOREclkx5,    	//PLL output on global n/w
  output [9:0] RAWDATAch0,     //Recovered ch 0 10-bit data 
  output [9:0] RAWDATAch1,     //Recovered ch 1 10-bit data
  output [9:0] RAWDATAch2,      //Recovered ch 2 10-bit data
  input	EXTFEEDBACK,  			//Driven by core logic. Not required HDMI mode.
  input	[7:0] DYNAMICDELAY,  	//Driven by core logic. Not required for HDMI mode.
  input	BYPASS,				//Driven by core logic. Not required for HDMI mode.
  input	LATCHINPUTVALUE, 	//iCEGate signal. Not required for HDMI mode
//Test Pins
  output	SDO,				//Output of PLL
  input	SDI,				//Driven by core logic
  input	SCLK				//Driven by core logic
  );

parameter FEEDBACK_PATH = "PHASE_AND_DELAY";	
parameter DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED"; 
parameter DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED"; 
parameter SHIFTREG_DIV_MODE = 2'b11; 	//Divide by 5.
parameter FDA_FEEDBACK = 4'b0000; 		//Integer 
parameter FDA_RELATIVE = 4'b0000; 		//Integer 
parameter PLLOUT_SELECT_PORTA = "GENCLK"; // Clkx5
parameter PLLOUT_SELECT_PORTB = "SHIFTREG_0deg"; // Clkx1

//Frequency Parameters: Current defaults are for TMDS Clk = 30-40MHz
parameter DIVR = 4'b0000; 	
parameter DIVF = 7'b0000000; 		// 7'b0000100; 
parameter DIVQ = 3'b010; 	
parameter FILTER_RANGE = 3'b011; 	

//Additional cbits
parameter ENABLE_ICEGATE_PORTA = 1'b0;
parameter ENABLE_ICEGATE_PORTB = 1'b0;

//Test Mode parameter
parameter TEST_MODE = 1'b0;
parameter EXTERNAL_DIVIDE_FACTOR = 1; //Not used by model. Added for PLL Config GUI.


    	wire clk1xout_global, clk5xout_global;  
    	wire clk1xout_core, clk5xout_core; 
  
  	wire ch0_clk5xin; 
  	wire ch1_clk5xin; 
  	wire ch2_clk5xin; 					
  
  SB_PLL40_2F_PAD_DS  dviphyPLL_i (
		.PACKAGEPIN(TMDSclkp),		
		.PACKAGEPINB(TMDSclkn),		
		.PLLOUTCOREA(clk5xout_core),		
		.PLLOUTGLOBALA(clk5xout_global),	
       		.PLLOUTCOREB(clk1xout_core),	
		.PLLOUTGLOBALB(clk1xout_global),	
		.EXTFEEDBACK(),  		
		.DYNAMICDELAY(),	
		.LOCK(PLLlock),			
		.BYPASS(1'b0),				
		.RESETB(RSTNpll),				
		.SDI(SDI),				
		.SDO(SDO),				
		.SCLK(SCLK),			
		.LATCHINPUTVALUE(1'b0)
	);

	defparam dviphyPLL_i.FEEDBACK_PATH = FEEDBACK_PATH ;   
	defparam dviphyPLL_i.DELAY_ADJUSTMENT_MODE_FEEDBACK = DELAY_ADJUSTMENT_MODE_FEEDBACK ; 
	defparam dviphyPLL_i.DELAY_ADJUSTMENT_MODE_RELATIVE = DELAY_ADJUSTMENT_MODE_RELATIVE ; 
	defparam dviphyPLL_i.SHIFTREG_DIV_MODE = SHIFTREG_DIV_MODE ; 
	defparam dviphyPLL_i.FDA_FEEDBACK = FDA_FEEDBACK ; 
	defparam dviphyPLL_i.FDA_RELATIVE = FDA_RELATIVE ;  
	defparam dviphyPLL_i.PLLOUT_SELECT_PORTA = PLLOUT_SELECT_PORTA ; 
	defparam dviphyPLL_i.PLLOUT_SELECT_PORTB = PLLOUT_SELECT_PORTB ; 
	defparam dviphyPLL_i.DIVR = DIVR ; 
	defparam dviphyPLL_i.DIVF = DIVF ; 
	defparam dviphyPLL_i.DIVQ = DIVQ ; 
	defparam dviphyPLL_i.FILTER_RANGE  = FILTER_RANGE ; 
	defparam dviphyPLL_i.ENABLE_ICEGATE_PORTA = ENABLE_ICEGATE_PORTA ; 
	defparam dviphyPLL_i.ENABLE_ICEGATE_PORTB = ENABLE_ICEGATE_PORTB ; 
	defparam dviphyPLL_i.TEST_MODE = TEST_MODE ; 
	defparam dviphyPLL_i.EXTERNAL_DIVIDE_FACTOR = EXTERNAL_DIVIDE_FACTOR ; 
	
	
	assign PLLOUTGLOBALclkx1 =  clk1xout_global ;  
	assign PLLOUTCOREclkx1   =  clk1xout_core; 
	assign PLLOUTGLOBALclkx5 =  clk5xout_global; 
	assign PLLOUTCOREclkx5   =  clk5xout_core; 
	
	//  -- channel 0  	
	clkdelay16  clkdelay16_ch0_i (
		.dlyin(clk5xout_global), 
		.dlyout(ch0_clk5xin), 
		.dly_sel(PHASELch0) 
	);
	
	dvi_deserializer deserializer_ch0_i (
		.en(EN),							
		.rstn(RSTNdeser), 	 
		.din(TMDSch0p), 
		.clkx5in(ch0_clk5xin),	
		.clkx1in(TMDSclkp),
		.rawdata(RAWDATAch0) 
	); 
	// -- channel 1 	
	clkdelay16  clkdelay16_ch1_i (
		.dlyin(clk5xout_global), 
		.dlyout(ch1_clk5xin), 
		.dly_sel(PHASELch1) 
	);								
	
	dvi_deserializer deserializer_ch1_i (
		.en(EN),							
		.rstn(RSTNdeser), 	 
		.din(TMDSch1p), 
		.clkx5in(ch1_clk5xin),	
		.clkx1in(TMDSclkp),
		.rawdata(RAWDATAch1) 
	); 
	
	// -- Channel 2 
	clkdelay16  clkdelay16_ch2_i (
		.dlyin(clk5xout_global), 
		.dlyout(ch2_clk5xin), 
		.dly_sel(PHASELch2) 
	);
	
	dvi_deserializer deserializer_ch2_i (
		.en(EN),							
		.rstn(RSTNdeser), 	 
		.din(TMDSch2p), 
		.clkx5in(ch2_clk5xin),	
		.clkx1in(TMDSclkp),
		.rawdata(RAWDATAch2) 
	); 


`ifdef TIMINGCHECK
specify
    // tp & tCQ arcs 
   (TMDSclkp *> PLLOUTGLOBALclkx1 ) = (1.0, 1.0);
   (TMDSclkp *> PLLOUTCOREclkx1 ) = (1.0, 1.0);	
   (TMDSclkp *> PLLOUTGLOBALclkx5  ) = (1.0, 1.0);	  
   (TMDSclkp *> PLLOUTCOREclkx5  ) = (1.0, 1.0); 

   (TMDSclkp *> RAWDATAch0[0]) = (1.0, 1.0);	
   (TMDSclkp *> RAWDATAch0[1]) = (1.0, 1.0);	
   (TMDSclkp *> RAWDATAch0[2]) = (1.0, 1.0);	
   (TMDSclkp *> RAWDATAch0[3]) = (1.0, 1.0);	
   (TMDSclkp *> RAWDATAch0[4]) = (1.0, 1.0);	
   (TMDSclkp *> RAWDATAch0[5]) = (1.0, 1.0);	
   (TMDSclkp *> RAWDATAch0[6]) = (1.0, 1.0);	
   (TMDSclkp *> RAWDATAch0[7]) = (1.0, 1.0);	
   (TMDSclkp *> RAWDATAch0[8]) = (1.0, 1.0);	 
   (TMDSclkp *> RAWDATAch0[9]) = (1.0, 1.0);	 

   (TMDSclkp *> RAWDATAch1[0]) = (1.0, 1.0);	
   (TMDSclkp *> RAWDATAch1[1]) = (1.0, 1.0);	
   (TMDSclkp *> RAWDATAch1[2]) = (1.0, 1.0);	
   (TMDSclkp *> RAWDATAch1[3]) = (1.0, 1.0);	
   (TMDSclkp *> RAWDATAch1[4]) = (1.0, 1.0);	
   (TMDSclkp *> RAWDATAch1[5]) = (1.0, 1.0);	
   (TMDSclkp *> RAWDATAch1[6]) = (1.0, 1.0);	
   (TMDSclkp *> RAWDATAch1[7]) = (1.0, 1.0);	
   (TMDSclkp *> RAWDATAch1[8]) = (1.0, 1.0);	 
   (TMDSclkp *> RAWDATAch1[9]) = (1.0, 1.0);	 

   (TMDSclkp *> RAWDATAch2[0]) = (1.0, 1.0);	
   (TMDSclkp *> RAWDATAch2[1]) = (1.0, 1.0);	
   (TMDSclkp *> RAWDATAch2[2]) = (1.0, 1.0);	
   (TMDSclkp *> RAWDATAch2[3]) = (1.0, 1.0);	
   (TMDSclkp *> RAWDATAch2[4]) = (1.0, 1.0);	
   (TMDSclkp *> RAWDATAch2[5]) = (1.0, 1.0);	
   (TMDSclkp *> RAWDATAch2[6]) = (1.0, 1.0);	
   (TMDSclkp *> RAWDATAch2[7]) = (1.0, 1.0);	
   (TMDSclkp *> RAWDATAch2[8]) = (1.0, 1.0);	 
   (TMDSclkp *> RAWDATAch2[9]) = (1.0, 1.0);	 


   // channel 0 setup-hold cheks 
   $setup(posedge TMDSch0p, posedge TMDSclkp, 1.0);
   $setup(negedge TMDSch0p, posedge TMDSclkp, 1.0);
   $hold (posedge TMDSclkp, posedge TMDSch0p, 1.0);
   $hold (posedge TMDSclkp, negedge TMDSch0p, 1.0);   
   $setup(posedge TMDSch0p, negedge TMDSclkp, 1.0);
   $setup(negedge TMDSch0p, negedge TMDSclkp, 1.0);
   $hold (negedge TMDSclkp, posedge TMDSch0p, 1.0);
   $hold (negedge TMDSclkp, negedge TMDSch0p, 1.0);
   
   $setup(posedge TMDSch0n, posedge TMDSclkp, 1.0);
   $setup(negedge TMDSch0n, posedge TMDSclkp, 1.0);
   $hold (posedge TMDSclkp, posedge TMDSch0n, 1.0);
   $hold (posedge TMDSclkp, negedge TMDSch0n, 1.0);   
   $setup(posedge TMDSch0n, negedge TMDSclkp, 1.0);
   $setup(negedge TMDSch0n, negedge TMDSclkp, 1.0);
   $hold (negedge TMDSclkp, posedge TMDSch0n, 1.0);
   $hold (negedge TMDSclkp, negedge TMDSch0n, 1.0);
	
   // channel 1 setup-hold cheks 
   $setup(posedge TMDSch1p, posedge TMDSclkp, 1.0);
   $setup(negedge TMDSch1p, posedge TMDSclkp, 1.0);
   $hold (posedge TMDSclkp, posedge TMDSch1p, 1.0);
   $hold (posedge TMDSclkp, negedge TMDSch1p, 1.0);   
   $setup(posedge TMDSch1p, negedge TMDSclkp, 1.0);
   $setup(negedge TMDSch1p, negedge TMDSclkp, 1.0);
   $hold (negedge TMDSclkp, posedge TMDSch1p, 1.0);
   $hold (negedge TMDSclkp, negedge TMDSch1p, 1.0);
   
   $setup(posedge TMDSch1n, posedge TMDSclkp, 1.0);
   $setup(negedge TMDSch1n, posedge TMDSclkp, 1.0);
   $hold (posedge TMDSclkp, posedge TMDSch1n, 1.0);
   $hold (posedge TMDSclkp, negedge TMDSch1n, 1.0);   
   $setup(posedge TMDSch1n, negedge TMDSclkp, 1.0);
   $setup(negedge TMDSch1n, negedge TMDSclkp, 1.0);
   $hold (negedge TMDSclkp, posedge TMDSch1n, 1.0);
   $hold (negedge TMDSclkp, negedge TMDSch1n, 1.0);


   // channel 2 setup-hold cheks 
   $setup(posedge TMDSch2p, posedge TMDSclkp, 1.0);
   $setup(negedge TMDSch2p, posedge TMDSclkp, 1.0);
   $hold (posedge TMDSclkp, posedge TMDSch2p, 1.0);
   $hold (posedge TMDSclkp, negedge TMDSch2p, 1.0);   
   $setup(posedge TMDSch2p, negedge TMDSclkp, 1.0);
   $setup(negedge TMDSch2p, negedge TMDSclkp, 1.0);
   $hold (negedge TMDSclkp, posedge TMDSch2p, 1.0);
   $hold (negedge TMDSclkp, negedge TMDSch2p, 1.0);
   
   $setup(posedge TMDSch2n, posedge TMDSclkp, 1.0);
   $setup(negedge TMDSch2n, posedge TMDSclkp, 1.0);
   $hold (posedge TMDSclkp, posedge TMDSch2n, 1.0);
   $hold (posedge TMDSclkp, negedge TMDSch2n, 1.0);   
   $setup(posedge TMDSch2n, negedge TMDSclkp, 1.0);
   $setup(negedge TMDSch2n, negedge TMDSclkp, 1.0);
   $hold (negedge TMDSclkp, posedge TMDSch2n, 1.0);
   $hold (negedge TMDSclkp, negedge TMDSch2n, 1.0);

endspecify
`endif   

	
endmodule  


//---------------------------------------//
//-------- 16 tap delay logic -----------//
//---------------------------------------//

`timescale 1ps /1ps 

module  clkdelay16 (
		dlyin, 
		dlyout, 
		dly_sel 
	);

parameter BUF_DELAY=100;	  	// 100ps +-25 ps 

input 			dlyin;  	// data to delay tap 
input 	[3:0]  		dly_sel;	// dealy adjustment. 0 - Nodelay    
output 			dlyout;      	// Delayed Data Line output   

wire 	[15:0] 	buf_y; 
reg         	delayed_data; 

// 16 tap buffer
assign  		 buf_y[0] = dlyin ; 	   
buf #BUF_DELAY  bufinst1 (buf_y[1],buf_y[0]);   
buf #BUF_DELAY  bufinst2 (buf_y[2],buf_y[1]);   
buf #BUF_DELAY  bufinst3 (buf_y[3],buf_y[2]);   
buf #BUF_DELAY  bufinst4 (buf_y[4],buf_y[3]);   
buf #BUF_DELAY  bufinst5 (buf_y[5],buf_y[4]);   
buf #BUF_DELAY  bufinst6 (buf_y[6],buf_y[5]);   
buf #BUF_DELAY  bufinst7 (buf_y[7],buf_y[6]);   
buf #BUF_DELAY  bufinst8 (buf_y[8],buf_y[7]);   
buf #BUF_DELAY  bufinst9 (buf_y[9],buf_y[8]);   
buf #BUF_DELAY  bufinst10 (buf_y[10],buf_y[9]); 
buf #BUF_DELAY  bufinst11 (buf_y[11],buf_y[10]);
buf #BUF_DELAY  bufinst12 (buf_y[12],buf_y[11]);
buf #BUF_DELAY  bufinst13 (buf_y[13],buf_y[12]);
buf #BUF_DELAY  bufinst14 (buf_y[14],buf_y[13]);
buf #BUF_DELAY  bufinst15 (buf_y[15],buf_y[14]);

// delay_sel mux 
always @*
begin 
	case(dly_sel) 
	4'd0: delayed_data  = buf_y[0];   
	4'd1: delayed_data  = buf_y[1];    
	4'd2: delayed_data  = buf_y[2];  
	4'd3: delayed_data  = buf_y[3];
	4'd4: delayed_data  = buf_y[4];
	4'd5: delayed_data  = buf_y[5];
	4'd6: delayed_data  = buf_y[6];
	4'd7: delayed_data  = buf_y[7];
	4'd8: delayed_data  = buf_y[8];
	4'd9: delayed_data  = buf_y[9];
	4'd10: delayed_data = buf_y[10];
	4'd11: delayed_data = buf_y[11];
	4'd12: delayed_data = buf_y[12];
	4'd13: delayed_data = buf_y[13];
	4'd14: delayed_data = buf_y[14];
	4'd15: delayed_data = buf_y[15];
	endcase
end 

assign dlyout = delayed_data ; 

endmodule

///--------------------------------------------------------------//
///----              dvi_deserializer			 -------//
///-------------------------------------------------------------// 

`timescale 1ns /1ps 
module dvi_deserializer (
	en,							
	rstn, 	 
	din, 
	clkx5in,	
	clkx1in,
	rawdata 
	); 

///---------------------------------------------------------/// 		
output reg  [9:0] rawdata ;		  // 10 bit raw data output 
input  rstn ;					  // Active low  deserializer reset 						  	
input  clkx5in ;				  // 5x clk input 
input  din ;					  // input stream 
input  clkx1in ;				 // 1x clk input 
input  en ;						 // global - clock enable 
///-----------------------------------------------------------///
wire 		clkx1 , clkx5 ; 
reg  		din_n0, din_n1;
reg 		din_p0; 
reg	[9:0] 	datain; 
wire [9:0]  mem_rdout;

assign 	clkx1 = clkx1in & en ; 
assign 	clkx5 = clkx5in & en ; 

/// ------------ Data Sampling Section  --------------- 
always@(negedge clkx5) 
begin
   if(en == 1'b1) 
	din_n0 <= din; 
end 

always@(posedge clkx5) 
begin 
	din_n1    <= ~din_n0;
	datain[8] <= din_n1; 
	datain[6] <= datain[8]; 
	datain[4] <= datain[6]; 
	datain[2] <= datain[4]; 
	datain[0] <= datain[2]; 
end 

always@(posedge clkx5) 
begin 
	din_p0 <= din; 
end 

always@(posedge clkx5) 
begin 
	datain[9] <= ~din_p0; 
	datain[7] <= datain[9]; 	
	datain[5] <= datain[7]; 
	datain[3] <= datain[5]; 
	datain[1] <= datain[3]; 
end 
	
reg [9:0]  datain_q;

always@(posedge clkx5) 	  
	begin 
	datain_q<=datain; 
end 
	
  reg 	[2:0]  	n_state; 
  reg 	[2:0]	p_state; 


  parameter ST0 = 3'b000;
  parameter ST1 = 3'b001;
  parameter ST2 = 3'b010;
  parameter ST3 = 3'b011;
  parameter ST4 = 3'b100;
  
  
  always@(p_state or rstn ) 
  begin 
	  case(p_state)
		  ST0 : begin  
		  		if (rstn==1'b1) n_state <= ST1; else n_state <= ST0;
		  		end  
		  ST1 : begin  
		  		if (rstn==1'b1) n_state <= ST2; else n_state <= ST1;
		  		end  	   
		  
		  ST2 : begin  
		  		if (rstn==1'b1) n_state <= ST3; else n_state <= ST2;
		  		end  
		  ST3 : begin  
		  		if (rstn==1'b1) n_state <= ST4; else n_state <= ST2;
		  		end  
		  default: n_state <=ST0; 
	  endcase
  end 
  
  always@(posedge clkx5 or negedge rstn) 
  begin 
	  if(rstn == 1'b0) 
		  p_state <= ST0; 
	  else if(en ==1'b1)
		  p_state <= n_state; 
 end 
 
 wire pulse_5cnt;
 reg sync_wren;
 
 assign pulse_5cnt = (p_state == ST3);	  
 
 always@(posedge clkx5) 
 begin 
	sync_wren <= pulse_5cnt;  
 end 
 				   
 // syncronous read , write reset signal gen 
  reg  rstsync_w, rstsync_r , wa_rst , ra_rst;						
  
  always@(posedge clkx5)
  begin 
	  rstsync_w <= rstn; 
	  rstsync_r <= rstsync_w; 
	  wa_rst    <= rstsync_r;				 
  //	  ra_rst 	<= wa_rst; 
  end 
 

  reg [3:0]  sync_rden; 

  
  always@(posedge clkx5)  // delay ra_rst 
  begin 
	sync_rden[0] <= rstsync_r;   
  	sync_rden[1] <= sync_rden[0];
	sync_rden[2] <= sync_rden[1];
	sync_rden[3] <= sync_rden[2];
	ra_rst <= sync_rden[3]; 
  end 
 
  //Address Generation Logics 
  reg [1:0] wa; 
  reg [1:0] ra; 
  
  always@(posedge clkx5 or negedge wa_rst)
  begin 
	  if(wa_rst == 1'b0) 
		  wa <= 2'b0;
	else if (sync_wren == 1'b1) 
		wa <= wa +1 ;     
  end 
		
  always @(posedge clkx1 or negedge ra_rst )
  begin 								   
	  if(ra_rst == 1'b0) 
		  ra <= 2'b0; 
	  else 
  	 	ra <= ra +1;  
  end  	    
  
  mem4x10  mem4x10_i 
  (
  .WDATAIN(datain_q),
  .WCLK(clkx5),
  .WE(sync_wren),
  .WADDR(wa),
  .RADDR(ra), 
  .RDATAOUT(mem_rdout)
  ); 
  
 always @ (posedge clkx1) begin
    rawdata<=mem_rdout;
 end		  
  
endmodule  

`timescale 1ns/1ps 
module mem4x10 (WDATAIN,WCLK,WE,WADDR,RADDR, RDATAOUT); 
	input [9:0]  WDATAIN; 
	input WCLK; 
	input WE; 
	input [1:0] WADDR;
	input [1:0] RADDR; 
	output [9:0] RDATAOUT; 
	
	reg [9:0] mem[0:3]; 
	
	// read first memory 
	always@(posedge WCLK) 
    	begin 		
		if(WE ==1'b1) begin 
			mem[WADDR] <= WDATAIN; 			
		end 					
    	end 						  	
	assign RDATAOUT = mem[RADDR];     

endmodule 	 


`timescale 1ps/1ps	
module SB_PLL40_2F_PAD_DS (
		PACKAGEPIN,		
		PACKAGEPINB,		
		PLLOUTCOREA,		//DIN0 output to core logic
		PLLOUTGLOBALA,	   	//PLL output to global network
        PLLOUTCOREB,		//PLL output to core logic
		PLLOUTGLOBALB,	   	//PLL output to global network
		EXTFEEDBACK,  			//Driven by core logic
		DYNAMICDELAY,		//Driven by core logic
		LOCK,				//Output of PLL
		BYPASS,				//Driven by core logic
		RESETB,				//Driven by core logic
		SDI,				//Driven by core logic. Test Pin
		SDO,				//Output to RB Logic Tile. Test Pin
		SCLK,				//Driven by core logic. Test Pin
		LATCHINPUTVALUE 	//iCEGate signal
);
inout 	PACKAGEPIN;		
inout 	PACKAGEPINB;		
output  PLLOUTCOREA;		//PLL output to core logic
output	PLLOUTGLOBALA;	   	//PLL output to global network
output  PLLOUTCOREB;		//PLL output to core logic
output	PLLOUTGLOBALB;	   	//PLL output to global network
input	EXTFEEDBACK;  			//Driven by core logic
input	[7:0] DYNAMICDELAY;  	//Driven by core logic
output	LOCK;				//Output of PLL
input	BYPASS;				//Driven by core logic
input	RESETB;				//Driven by core logic
input	LATCHINPUTVALUE; 	//iCEGate signal
//Test Pins
output	SDO;				//Output of PLL
input	SDI;				//Driven by core logic
input	SCLK;				//Driven by core logic

//Feedback
parameter FEEDBACK_PATH = "SIMPLE";	//String  (simple, delay, phase_and_delay, external) 
parameter DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED"; 
parameter DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED"; 
parameter SHIFTREG_DIV_MODE = 2'b00; //00-->Divide by 4, 01-->Divide by 7, 11-->Divide by 5.
parameter FDA_FEEDBACK = 4'b0000; 		//Integer. 

//Output 
parameter FDA_RELATIVE = 4'b0000; 		//Integer. 
parameter PLLOUT_SELECT_PORTA = "GENCLK"; //
parameter PLLOUT_SELECT_PORTB = "GENCLK"; //

//Use the Spreadsheet to populate the values below.
parameter DIVR = 4'b0000; 	//determine a good default value
parameter DIVF = 7'b0000000; //determine a good default value
parameter DIVQ = 3'b000; 	//determine a good default value
parameter FILTER_RANGE = 3'b000; 	//determine a good default value

//Additional cbits
parameter ENABLE_ICEGATE_PORTA = 1'b0;
parameter ENABLE_ICEGATE_PORTB = 1'b0;

//Test Mode parameter
parameter TEST_MODE = 1'b0;
parameter EXTERNAL_DIVIDE_FACTOR = 1; //Not used by model. Added for PLL Config GUI.

wire SPLLOUT1net , SPLLOUT2net; 

SbtSPLL40 instSbtSPLL (
		.REFERENCECLK (PACKAGEPIN),
		.EXTFEEDBACK (EXTFEEDBACK),  	
		.DYNAMICDELAY (DYNAMICDELAY),		
		.BYPASS (BYPASS),
		.RESETB (~RESETB),	
		
		.PLLOUT1 (SPLLOUT1net),	
		.PLLOUT2 (SPLLOUT2net),		
		.LOCK (LOCK)   	

);
defparam instSbtSPLL.DIVR = DIVR;	
defparam instSbtSPLL.DIVF = DIVF;
defparam instSbtSPLL.DIVQ = DIVQ;
defparam instSbtSPLL.FILTER_RANGE = FILTER_RANGE;
defparam instSbtSPLL.FEEDBACK_PATH = FEEDBACK_PATH;
defparam instSbtSPLL.DELAY_ADJUSTMENT_MODE_RELATIVE = DELAY_ADJUSTMENT_MODE_RELATIVE;
defparam instSbtSPLL.DELAY_ADJUSTMENT_MODE_FEEDBACK = DELAY_ADJUSTMENT_MODE_FEEDBACK;
defparam instSbtSPLL.SHIFTREG_DIV_MODE = SHIFTREG_DIV_MODE;
defparam instSbtSPLL.FDA_RELATIVE = FDA_RELATIVE; 
defparam instSbtSPLL.FDA_FEEDBACK = FDA_FEEDBACK; 
defparam instSbtSPLL.PLLOUT_SELECT_PORTA = PLLOUT_SELECT_PORTA;
defparam instSbtSPLL.PLLOUT_SELECT_PORTB = PLLOUT_SELECT_PORTB;

assign PLLOUTCOREA = ((ENABLE_ICEGATE_PORTA != 0) && LATCHINPUTVALUE) ? PLLOUTCOREA : SPLLOUT1net;
assign PLLOUTGLOBALA = ((ENABLE_ICEGATE_PORTA != 0) && LATCHINPUTVALUE)  ? PLLOUTGLOBALA : SPLLOUT1net;
assign PLLOUTCOREB = ((ENABLE_ICEGATE_PORTB != 0) && LATCHINPUTVALUE) ? PLLOUTCOREB : SPLLOUT2net;
assign PLLOUTGLOBALB = ((ENABLE_ICEGATE_PORTB != 0) && LATCHINPUTVALUE)  ? PLLOUTGLOBALB : SPLLOUT2net;

`ifdef TIMINGCHECK
specify
   (PACKAGEPIN *> PLLOUTGLOBALA) = (1.0, 1.0);
   (PACKAGEPIN *> PLLOUTCOREA) = (1.0, 1.0);
   (PACKAGEPIN *> PLLOUTGLOBALB) = (1.0, 1.0);
   (PACKAGEPIN *> PLLOUTCOREB) = (1.0, 1.0);

endspecify
`endif

endmodule // SB_PLL40_2F_PAD_DS



`timescale 1ps/1ps
module SB_PLL40_PAD_DS (
		PACKAGEPIN,		
		PACKAGEPINB,		
		PLLOUTCORE,		//PLL output to core logic
		PLLOUTGLOBAL,	   	//PLL output to global network
		EXTFEEDBACK,  			//Driven by core logic
		DYNAMICDELAY,		//Driven by core logic
		LOCK,				//Output of PLL
		BYPASS,				//Driven by core logic
		RESETB,				//Driven by core logic
		SDI,				//Driven by core logic. Test Pin
		SDO,				//Output to RB Logic Tile. Test Pin
		SCLK,				//Driven by core logic. Test Pin
		LATCHINPUTVALUE 	//iCEGate signal
);
inout 	PACKAGEPIN;		
inout 	PACKAGEPINB;		
output 	PLLOUTCORE;		//PLL output to core logic
output	PLLOUTGLOBAL;	   	//PLL output to global network
input	EXTFEEDBACK;  			//Driven by core logic
input	[7:0] DYNAMICDELAY;  	//Driven by core logic
output	LOCK;				//Output of PLL
input	BYPASS;				//Driven by core logic
input	RESETB;				//Driven by core logic
input	LATCHINPUTVALUE; 	//iCEGate signal
//Test Pins
output	SDO;				//Output of PLL
input	SDI;				//Driven by core logic
input	SCLK;				//Driven by core logic


//Feedback
parameter FEEDBACK_PATH = "SIMPLE";	//String  (simple, delay, phase_and_delay, external) 
parameter DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED"; 
parameter DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED"; 
parameter SHIFTREG_DIV_MODE = 2'b00; //00-->Divide by 4, 01-->Divide by 7, 11-->Divide by 5.
parameter FDA_FEEDBACK = 4'b0000; 		//Integer. 

parameter FDA_RELATIVE = 4'b0000; 		//Integer. 
parameter PLLOUT_SELECT = "GENCLK"; //

//Use the Spreadsheet to populate the values below.
parameter DIVR = 4'b0000; 	//determine a good default value
parameter DIVF = 7'b0000000; //determine a good default value
parameter DIVQ = 3'b000; 	//determine a good default value
parameter FILTER_RANGE = 3'b000; 	//determine a good default value

//Additional cbits
parameter ENABLE_ICEGATE = 1'b0;

//Test Mode parameter
parameter TEST_MODE = 1'b0;
parameter EXTERNAL_DIVIDE_FACTOR = 1; //Not used by model. Added for PLL Config GUI.

wire SPLLOUT1net,SPLLOUT2net; 

SbtSPLL40 instSbtSPLL (
		.REFERENCECLK (PACKAGEPIN),
		.EXTFEEDBACK (EXTFEEDBACK),  	
		.DYNAMICDELAY (DYNAMICDELAY),		
		.BYPASS (BYPASS),
		.RESETB (~RESETB),	
		
		.PLLOUT1 (SPLLOUT1net),	
		.PLLOUT2 (SPLLOUT2net),		
		.LOCK (LOCK)   	

);
defparam instSbtSPLL.DIVR = DIVR;	
defparam instSbtSPLL.DIVF = DIVF;
defparam instSbtSPLL.DIVQ = DIVQ;
defparam instSbtSPLL.FILTER_RANGE = FILTER_RANGE;
defparam instSbtSPLL.FEEDBACK_PATH = FEEDBACK_PATH;
defparam instSbtSPLL.DELAY_ADJUSTMENT_MODE_RELATIVE = DELAY_ADJUSTMENT_MODE_RELATIVE;
defparam instSbtSPLL.DELAY_ADJUSTMENT_MODE_FEEDBACK = DELAY_ADJUSTMENT_MODE_FEEDBACK;
defparam instSbtSPLL.SHIFTREG_DIV_MODE = SHIFTREG_DIV_MODE;
defparam instSbtSPLL.FDA_RELATIVE = FDA_RELATIVE; 
defparam instSbtSPLL.FDA_FEEDBACK = FDA_FEEDBACK; 
defparam instSbtSPLL.PLLOUT_SELECT_PORTA = PLLOUT_SELECT;
defparam instSbtSPLL.PLLOUT_SELECT_PORTB = "GENCLK";


assign PLLOUTCORE = ((ENABLE_ICEGATE != 0) && LATCHINPUTVALUE) ? PLLOUTCORE : SPLLOUT1net;
assign PLLOUTGLOBAL = ((ENABLE_ICEGATE != 0) && LATCHINPUTVALUE)  ? PLLOUTGLOBAL : SPLLOUT1net;

`ifdef TIMINGCHECK
specify
   (PACKAGEPIN *> PLLOUTGLOBAL) = (1.0, 1.0);
   (PACKAGEPIN *> PLLOUTCORE) = (1.0, 1.0);
endspecify
`endif

endmodule // SB_PLL40_PAD_DS
 

//-----------------------------------------------// 
//----	SB_MAC16 DSP Primitive             ------//
//-----------------------------------------------// 
`timescale 1ps/1ps
module SB_MAC16 (
		A,
		B,
		C,
		D,
		O,
		CLK,
		CE,
		IRSTTOP,
	    IRSTBOT,
		ORSTTOP,
		ORSTBOT,
		AHOLD,
		BHOLD,
		CHOLD,
		DHOLD,
		OHOLDTOP,
		OHOLDBOT,
		OLOADTOP,
		OLOADBOT,
		ADDSUBTOP,
		ADDSUBBOT,
		CO,
		CI,  		//from bottom tile
		ACCUMCI, 	// Carry input from MAC CO below
		ACCUMCO, 	// Carry output to above MAC block.    
		SIGNEXTIN,
		SIGNEXTOUT
);
output 	[31:0] O;	 // Output [31:0]
input	[15:0] A;        // data  to upper mult block / upper accum block.
input	[15:0] B;        // data  to lower mult block / lower accum block.   
input	[15:0] C;        // direct data  to upper accum block. 
input	[15:0] D;        // direct data  to lower accum block.
input	CLK;	         // Clock for MAC16 elements 
input	CE;              // Clock enable . global control 
input	IRSTTOP;         // Active High  reset for  A,C registers,upper half multplier pipeline regs(16). 
input	IRSTBOT;         // Active High reset for  B,D registers, lower half multiplier pipeline regs(16), 32 bit result pipelines regs   
input	ORSTTOP;	 // Active High reset for top accum registers O[31:16]
input	ORSTBOT;         // Active High reset for bottom accum registers O[15:0]   
input   AHOLD;           // Active High hold data signal for A register
input   BHOLD;           // Active High hold data signal for B register   
input   CHOLD;           // Active High hold data signal for C register
input   DHOLD;           // Active High hold data signal for D register 
input   OHOLDTOP;        // Active High hold data signal for top accum registers O[31:16]
input   OHOLDBOT;        // Active High hold data signal for bottom  accum registers O[15:0]     
input 	OLOADTOP;        // Load top accum regiser with  direct input C or Registered data C.  
input 	OLOADBOT;        // Load bottom accum regisers with direct input D or Registered data D
input 	ADDSUBTOP;       // Control for Add/Sub operation for top accum . 0-addition , 1-subtraction.  
input 	ADDSUBBOT;       // Control for Add/Sub operation for bottom accum . 0-addition , 1-subtraction.
output  CO;              // top accumulator carry out to next LUT
input 	CI;              // bottom accumaltor carry in signal from lower LUT block. 
input   ACCUMCI;         // Carry in from  MAC16 below
output  ACCUMCO;         // Carry out to MAC16 above
input   SIGNEXTIN;	 // Single bit Sign extenstion from MAC16 below         
output  SIGNEXTOUT;      // Single bit Sign extenstion to MAC16 above


parameter NEG_TRIGGER = 1'b0;    
parameter C_REG = 1'b0;     			// C0
parameter A_REG = 1'b0;     			// C1
parameter B_REG = 1'b0;     			// C2
parameter D_REG = 1'b0;     			// C3

parameter TOP_8x8_MULT_REG = 1'b0; 		//C4
parameter BOT_8x8_MULT_REG = 1'b0; 		//C5
parameter PIPELINE_16x16_MULT_REG1 = 1'b0; 	//C6
parameter PIPELINE_16x16_MULT_REG2 = 1'b0; 	//C7

parameter TOPOUTPUT_SELECT =  2'b00; 		//COMB, ACCUM_REG, MULT_8x8, MULT_16x16  // {C9,C8} = 00, 01, 10, 11
parameter TOPADDSUB_LOWERINPUT = 2'b00; 	//DATA, MULT_8x8, MULT_16x16, SIGNEXT    // {C11,C10} = 00, 01, 10, 11
parameter TOPADDSUB_UPPERINPUT = 1'b0; 		//ACCUM_REG, DATAC  			 //  C12 = 0, 1
parameter TOPADDSUB_CARRYSELECT = 2'b00; 	//LOGIC0, LOGIC1, LCOCAS, GENERATED_CARRY (LCO) // {C14, C13} = 00, 01, 10, 11

parameter BOTOUTPUT_SELECT =  2'b00; 		//COMB, ACCUM_REG, MULT_8x8, MULT_16x16   // {C16,C15} = 00, 01, 10, 11
parameter BOTADDSUB_LOWERINPUT = 2'b00; 	//DATA, MULT_8x8, MULT_16x16, SIGNEXTIN   // {C18,C17} = 00, 01, 10, 11
parameter BOTADDSUB_UPPERINPUT = 1'b0;  	//ACCUM_REG, DATAD   			  // C19 = 0, 1
parameter BOTADDSUB_CARRYSELECT = 2'b00; 	//LOGIC0, LOGIC1, ACCUMCI, CI  		  // {C21, C20} = 00, 01, 10, 11
parameter MODE_8x8 = 1'b0; 			// C22 

parameter A_SIGNED = 1'b0;  			// C23
parameter B_SIGNED = 1'b0;  			// C24	 

//--------- local params ----------------------------------------------------// 
localparam cbits_inreg   	= {D_REG,B_REG,A_REG,C_REG}; 
localparam cbits_mpyreg   	= {PIPELINE_16x16_MULT_REG2,PIPELINE_16x16_MULT_REG1,BOT_8x8_MULT_REG,TOP_8x8_MULT_REG};
localparam cbits_topmac	 	= {TOPADDSUB_CARRYSELECT,TOPADDSUB_UPPERINPUT,TOPADDSUB_LOWERINPUT,TOPOUTPUT_SELECT};
localparam cbits_botmac	 	= {BOTADDSUB_CARRYSELECT,BOTADDSUB_UPPERINPUT,BOTADDSUB_LOWERINPUT,BOTOUTPUT_SELECT};
localparam cbits_sign	 	= {B_SIGNED,A_SIGNED,MODE_8x8}; 
localparam cbits 	  	= {cbits_sign,cbits_botmac,cbits_topmac,cbits_mpyreg,cbits_inreg}; 

wire CLK_g , intCLK; 
reg NOTIFIER;


//------------------- initial block --------------------------------------// 
	
	initial 
begin 
	
	
	
	if( (TOPOUTPUT_SELECT != 2'b00 )&& (TOPOUTPUT_SELECT != 2'b01 ) && (TOPOUTPUT_SELECT != 2'b10 ) && (TOPOUTPUT_SELECT !=2'b11 ) ) begin 
	$display("Error: TOPOUTPUT_SELECT parameter is set to incorrect value. Exiting Simulation ...."); 
	$finish;	
	end 
	if( (TOPADDSUB_LOWERINPUT != 2'b00) && (TOPADDSUB_LOWERINPUT != 2'b01) && (TOPADDSUB_LOWERINPUT != 2'b10) && (TOPADDSUB_LOWERINPUT != 2'b11) ) begin 
	$display("Error: TOPADDSUB_LOWERINPUT parameter is set to incorrect value. Exiting Simulation ...."); 
	$finish; 
	end 
	if( (TOPADDSUB_UPPERINPUT != 1'b0 ) && (TOPADDSUB_UPPERINPUT != 1'b1) ) begin
	$display("Error: TOPADDSUB_UPPERINPUT parameter is set to incorrect value. Exiting Simulation ....");
        $finish;
        end
	if( (TOPADDSUB_CARRYSELECT != 2'b00 )&&(TOPADDSUB_CARRYSELECT != 2'b01) && (TOPADDSUB_CARRYSELECT != 2'b10) &&(TOPADDSUB_CARRYSELECT != 2'b11)) begin 
	$display("Error: TOPADDSUB_CARRYSELECT parameter is set to incorrect value. Exiting Simulation ....");
        $finish;
        end

	
	if( (BOTOUTPUT_SELECT != 2'b00 )&& (BOTOUTPUT_SELECT != 2'b01 ) && (BOTOUTPUT_SELECT != 2'b10 ) && (BOTOUTPUT_SELECT !=2'b11 ) ) begin 
	$display("Error: BOTOUTPUT_SELECT parameter is set to incorrect value. Exiting Simulation ...."); 
	$finish;	
	end 
	if( (BOTADDSUB_LOWERINPUT != 2'b00) && (BOTADDSUB_LOWERINPUT != 2'b01) && (BOTADDSUB_LOWERINPUT != 2'b10) && (BOTADDSUB_LOWERINPUT != 2'b11) ) begin 
	$display("Error: BOTADDSUB_LOWERINPUT parameter is set to incorrect value. Exiting Simulation ...."); 
	$finish; 
	end 
	if( (BOTADDSUB_UPPERINPUT != 1'b0 ) && (BOTADDSUB_UPPERINPUT != 1'b1) ) begin
	$display("Error:BOTADDSUB_UPPERINPUT parameter is set to incorrect value. Exiting Simulation ....");
        $finish;
        end
	if( (BOTADDSUB_CARRYSELECT != 2'b00 ) && (BOTADDSUB_CARRYSELECT != 2'b01) && (BOTADDSUB_CARRYSELECT != 2'b10) && (BOTADDSUB_CARRYSELECT != 2'b11)) begin 
	$display("Error: BOTADDSUB_CARRYSELECT parameter is set to incorrect value. Exiting Simulation ....");
        $finish;
        end
	
	//Validation for mode8x8.
		if (PIPELINE_16x16_MULT_REG1 == 1'b1 || PIPELINE_16x16_MULT_REG2 ==1'b1 ) begin   		
		$display ("**************  INFO  ***********************************"); 
		$display ("Info : To Reset 16x16 multiplier INTERNAL PIPELINE REGISTER assert both IRSTTOP and IRSTBOT signals") ;  
	        $display ("Info : To Reset 16x16 multiplier OUTPUT  REGISTER   assert IRSTBOT signal");  	
		$display ("**********************************************************"); 	
		end else if ( (PIPELINE_16x16_MULT_REG1 == 1'b1 || PIPELINE_16x16_MULT_REG2 ==1'b1) &&  MODE_8x8 == 1'b1) begin
		  
		$display ("***********  ERROR  ****************************************"); 
		$display ("Error : MODE_8x8 parameter is set to 1. To use 16x16 mulitplier internal and output registers it should be set to 0.Exiting Simulation ...."); 
		
		$display ("***************************************************************"); 	
		$finish; 
		end else if( (PIPELINE_16x16_MULT_REG1 == 1'b0 &&  PIPELINE_16x16_MULT_REG2 ==1'b0)  &&  MODE_8x8 == 1'b0 ) begin
                $display ("************ WARNING  **********************************************");
                $display ("Warning : When 16x16 multiplier PIPELINE REGISTERS are not used, set MODE_8x8 to 1(power save mode) ");
                $display ("*******************************************************************");
		end 


end	// initial  

//-------------------------- Default input signals -------------------------------------// 
assign (weak0,weak1) CE 	= 1'b1; 
assign (weak0,weak1) A  	= 16'b0; 
assign (weak0,weak1) B  	= 16'b0; 
assign (weak0,weak1) C  	= 16'b0; 
assign (weak0,weak1) D  	= 16'b0; 
assign (weak0,weak1) AHOLD 	= 1'b0; 
assign (weak0,weak1) BHOLD 	= 1'b0; 
assign (weak0,weak1) CHOLD 	= 1'b0; 
assign (weak0,weak1) DHOLD    	= 1'b0; 
assign (weak0,weak1) IRSTTOP  	= 1'b0; 
assign (weak0,weak1) IRSTBOT  	= 1'b0; 
assign (weak0,weak1) ORSTTOP  	= 1'b0; 
assign (weak0,weak1) ORSTBOT  	= 1'b0; 
assign (weak0,weak1) OLOADTOP 	= 1'b0; 
assign (weak0,weak1) OLOADBOT 	= 1'b0; 
assign (weak0,weak1) ADDSUBTOP	= 1'b0; 
assign (weak0,weak1) ADDSUBBOT  = 1'b0; 
assign (weak0,weak1) OHOLDTOP   = 1'b0; 
assign (weak0,weak1) OHOLDBOT	= 1'b0;   
assign (weak0,weak1) CI		= 1'b0;   
assign (weak0,weak1) ACCUMCI	= 1'b0;   


//---------------------------Logic section --------------------------------------------// 

assign CLK_g = (CLK & CE);  				// CE=0 disables entire clock  
assign intCLK = (CLK_g ^ NEG_TRIGGER);			// Clock Polarity control 

 mac16_physical  mac16physical_i (
	 .CLK(intCLK) ,
	 .A(A) ,
	 .B(B) ,
	 .C(C) ,
	 .D(D) ,
	 .IHRST(IRSTTOP),
	 .ILRST(IRSTBOT),
	 .OHRST(ORSTTOP),
	 .OLRST(ORSTBOT),
	 .AHLD(AHOLD),
	 .BHLD(BHOLD),
	 .CHLD(CHOLD),
	 .DHLD(DHOLD),
		
	 .OHHLD(OHOLDTOP),
	 .OLHLD(OHOLDBOT),
	 .OHADS(ADDSUBTOP),
	 .OLADS(ADDSUBBOT),
	 .OHLDA(OLOADTOP),
	 .OLLDA(OLOADBOT),
	 .CICAS(ACCUMCI),
	 .CI(CI),
	 .SIGNEXTIN(SIGNEXTIN),
	 .SIGNEXTOUT(SIGNEXTOUT),
	 .COCAS(ACCUMCO),
	 .CO(CO),
	 .O(O), 
	 .CBIT(cbits)
    );
`ifdef TIMINGCHECK		
specify


		 (A[0] *> O[0])=(0.0,0.0); 
        (A[0] *> O[1])=(0.0,0.0); 
        (A[0] *> O[2])=(0.0,0.0); 
        (A[0] *> O[3])=(0.0,0.0); 
        (A[0] *> O[4])=(0.0,0.0); 
        (A[0] *> O[5])=(0.0,0.0); 
        (A[0] *> O[6])=(0.0,0.0); 
        (A[0] *> O[7])=(0.0,0.0); 
        (A[0] *> O[8])=(0.0,0.0); 
        (A[0] *> O[9])=(0.0,0.0); 
        (A[0] *> O[10])=(0.0,0.0); 
        (A[0] *> O[11])=(0.0,0.0); 
        (A[0] *> O[12])=(0.0,0.0); 
        (A[0] *> O[13])=(0.0,0.0); 
        (A[0] *> O[14])=(0.0,0.0); 
        (A[0] *> O[15])=(0.0,0.0); 
        (A[0] *> O[16])=(0.0,0.0); 
        (A[0] *> O[17])=(0.0,0.0); 
        (A[0] *> O[18])=(0.0,0.0); 
        (A[0] *> O[19])=(0.0,0.0); 
        (A[0] *> O[20])=(0.0,0.0); 
        (A[0] *> O[21])=(0.0,0.0); 
        (A[0] *> O[22])=(0.0,0.0); 
        (A[0] *> O[23])=(0.0,0.0); 
        (A[0] *> O[24])=(0.0,0.0); 
        (A[0] *> O[25])=(0.0,0.0); 
        (A[0] *> O[26])=(0.0,0.0); 
        (A[0] *> O[27])=(0.0,0.0); 
        (A[0] *> O[28])=(0.0,0.0); 
        (A[0] *> O[29])=(0.0,0.0); 
        (A[0] *> O[30])=(0.0,0.0); 
        (A[0] *> O[31])=(0.0,0.0); 
        (A[1] *> O[0])=(0.0,0.0); 
        (A[1] *> O[1])=(0.0,0.0); 
        (A[1] *> O[2])=(0.0,0.0); 
        (A[1] *> O[3])=(0.0,0.0); 
        (A[1] *> O[4])=(0.0,0.0); 
        (A[1] *> O[5])=(0.0,0.0); 
        (A[1] *> O[6])=(0.0,0.0); 
        (A[1] *> O[7])=(0.0,0.0); 
        (A[1] *> O[8])=(0.0,0.0); 
        (A[1] *> O[9])=(0.0,0.0); 
        (A[1] *> O[10])=(0.0,0.0); 
        (A[1] *> O[11])=(0.0,0.0); 
        (A[1] *> O[12])=(0.0,0.0); 
        (A[1] *> O[13])=(0.0,0.0); 
        (A[1] *> O[14])=(0.0,0.0); 
        (A[1] *> O[15])=(0.0,0.0); 
        (A[1] *> O[16])=(0.0,0.0); 
        (A[1] *> O[17])=(0.0,0.0); 
        (A[1] *> O[18])=(0.0,0.0); 
        (A[1] *> O[19])=(0.0,0.0); 
        (A[1] *> O[20])=(0.0,0.0); 
        (A[1] *> O[21])=(0.0,0.0); 
        (A[1] *> O[22])=(0.0,0.0); 
        (A[1] *> O[23])=(0.0,0.0); 
        (A[1] *> O[24])=(0.0,0.0); 
        (A[1] *> O[25])=(0.0,0.0); 
        (A[1] *> O[26])=(0.0,0.0); 
        (A[1] *> O[27])=(0.0,0.0); 
        (A[1] *> O[28])=(0.0,0.0); 
        (A[1] *> O[29])=(0.0,0.0); 
        (A[1] *> O[30])=(0.0,0.0); 
        (A[1] *> O[31])=(0.0,0.0); 
        (A[2] *> O[0])=(0.0,0.0); 
        (A[2] *> O[1])=(0.0,0.0); 
        (A[2] *> O[2])=(0.0,0.0); 
        (A[2] *> O[3])=(0.0,0.0); 
        (A[2] *> O[4])=(0.0,0.0); 
        (A[2] *> O[5])=(0.0,0.0); 
        (A[2] *> O[6])=(0.0,0.0); 
        (A[2] *> O[7])=(0.0,0.0); 
        (A[2] *> O[8])=(0.0,0.0); 
        (A[2] *> O[9])=(0.0,0.0); 
        (A[2] *> O[10])=(0.0,0.0); 
        (A[2] *> O[11])=(0.0,0.0); 
        (A[2] *> O[12])=(0.0,0.0); 
        (A[2] *> O[13])=(0.0,0.0); 
        (A[2] *> O[14])=(0.0,0.0); 
        (A[2] *> O[15])=(0.0,0.0); 
        (A[2] *> O[16])=(0.0,0.0); 
        (A[2] *> O[17])=(0.0,0.0); 
        (A[2] *> O[18])=(0.0,0.0); 
        (A[2] *> O[19])=(0.0,0.0); 
        (A[2] *> O[20])=(0.0,0.0); 
        (A[2] *> O[21])=(0.0,0.0); 
        (A[2] *> O[22])=(0.0,0.0); 
        (A[2] *> O[23])=(0.0,0.0); 
        (A[2] *> O[24])=(0.0,0.0); 
        (A[2] *> O[25])=(0.0,0.0); 
        (A[2] *> O[26])=(0.0,0.0); 
        (A[2] *> O[27])=(0.0,0.0); 
        (A[2] *> O[28])=(0.0,0.0); 
        (A[2] *> O[29])=(0.0,0.0); 
        (A[2] *> O[30])=(0.0,0.0); 
        (A[2] *> O[31])=(0.0,0.0); 
        (A[3] *> O[0])=(0.0,0.0); 
        (A[3] *> O[1])=(0.0,0.0); 
        (A[3] *> O[2])=(0.0,0.0); 
        (A[3] *> O[3])=(0.0,0.0); 
        (A[3] *> O[4])=(0.0,0.0); 
        (A[3] *> O[5])=(0.0,0.0); 
        (A[3] *> O[6])=(0.0,0.0); 
        (A[3] *> O[7])=(0.0,0.0); 
        (A[3] *> O[8])=(0.0,0.0); 
        (A[3] *> O[9])=(0.0,0.0); 
        (A[3] *> O[10])=(0.0,0.0); 
        (A[3] *> O[11])=(0.0,0.0); 
        (A[3] *> O[12])=(0.0,0.0); 
        (A[3] *> O[13])=(0.0,0.0); 
        (A[3] *> O[14])=(0.0,0.0); 
        (A[3] *> O[15])=(0.0,0.0); 
        (A[3] *> O[16])=(0.0,0.0); 
        (A[3] *> O[17])=(0.0,0.0); 
        (A[3] *> O[18])=(0.0,0.0); 
        (A[3] *> O[19])=(0.0,0.0); 
        (A[3] *> O[20])=(0.0,0.0); 
        (A[3] *> O[21])=(0.0,0.0); 
        (A[3] *> O[22])=(0.0,0.0); 
        (A[3] *> O[23])=(0.0,0.0); 
        (A[3] *> O[24])=(0.0,0.0); 
        (A[3] *> O[25])=(0.0,0.0); 
        (A[3] *> O[26])=(0.0,0.0); 
        (A[3] *> O[27])=(0.0,0.0); 
        (A[3] *> O[28])=(0.0,0.0); 
        (A[3] *> O[29])=(0.0,0.0); 
        (A[3] *> O[30])=(0.0,0.0); 
        (A[3] *> O[31])=(0.0,0.0); 
        (A[4] *> O[0])=(0.0,0.0); 
        (A[4] *> O[1])=(0.0,0.0); 
        (A[4] *> O[2])=(0.0,0.0); 
        (A[4] *> O[3])=(0.0,0.0); 
        (A[4] *> O[4])=(0.0,0.0); 
        (A[4] *> O[5])=(0.0,0.0); 
        (A[4] *> O[6])=(0.0,0.0); 
        (A[4] *> O[7])=(0.0,0.0); 
        (A[4] *> O[8])=(0.0,0.0); 
        (A[4] *> O[9])=(0.0,0.0); 
        (A[4] *> O[10])=(0.0,0.0); 
        (A[4] *> O[11])=(0.0,0.0); 
        (A[4] *> O[12])=(0.0,0.0); 
        (A[4] *> O[13])=(0.0,0.0); 
        (A[4] *> O[14])=(0.0,0.0); 
        (A[4] *> O[15])=(0.0,0.0); 
        (A[4] *> O[16])=(0.0,0.0); 
        (A[4] *> O[17])=(0.0,0.0); 
        (A[4] *> O[18])=(0.0,0.0); 
        (A[4] *> O[19])=(0.0,0.0); 
        (A[4] *> O[20])=(0.0,0.0); 
        (A[4] *> O[21])=(0.0,0.0); 
        (A[4] *> O[22])=(0.0,0.0); 
        (A[4] *> O[23])=(0.0,0.0); 
        (A[4] *> O[24])=(0.0,0.0); 
        (A[4] *> O[25])=(0.0,0.0); 
        (A[4] *> O[26])=(0.0,0.0); 
        (A[4] *> O[27])=(0.0,0.0); 
        (A[4] *> O[28])=(0.0,0.0); 
        (A[4] *> O[29])=(0.0,0.0); 
        (A[4] *> O[30])=(0.0,0.0); 
        (A[4] *> O[31])=(0.0,0.0); 
        (A[5] *> O[0])=(0.0,0.0); 
        (A[5] *> O[1])=(0.0,0.0); 
        (A[5] *> O[2])=(0.0,0.0); 
        (A[5] *> O[3])=(0.0,0.0); 
        (A[5] *> O[4])=(0.0,0.0); 
        (A[5] *> O[5])=(0.0,0.0); 
        (A[5] *> O[6])=(0.0,0.0); 
        (A[5] *> O[7])=(0.0,0.0); 
        (A[5] *> O[8])=(0.0,0.0); 
        (A[5] *> O[9])=(0.0,0.0); 
        (A[5] *> O[10])=(0.0,0.0); 
        (A[5] *> O[11])=(0.0,0.0); 
        (A[5] *> O[12])=(0.0,0.0); 
        (A[5] *> O[13])=(0.0,0.0); 
        (A[5] *> O[14])=(0.0,0.0); 
        (A[5] *> O[15])=(0.0,0.0); 
        (A[5] *> O[16])=(0.0,0.0); 
        (A[5] *> O[17])=(0.0,0.0); 
        (A[5] *> O[18])=(0.0,0.0); 
        (A[5] *> O[19])=(0.0,0.0); 
        (A[5] *> O[20])=(0.0,0.0); 
        (A[5] *> O[21])=(0.0,0.0); 
        (A[5] *> O[22])=(0.0,0.0); 
        (A[5] *> O[23])=(0.0,0.0); 
        (A[5] *> O[24])=(0.0,0.0); 
        (A[5] *> O[25])=(0.0,0.0); 
        (A[5] *> O[26])=(0.0,0.0); 
        (A[5] *> O[27])=(0.0,0.0); 
        (A[5] *> O[28])=(0.0,0.0); 
        (A[5] *> O[29])=(0.0,0.0); 
        (A[5] *> O[30])=(0.0,0.0); 
        (A[5] *> O[31])=(0.0,0.0); 
        (A[6] *> O[0])=(0.0,0.0); 
        (A[6] *> O[1])=(0.0,0.0); 
        (A[6] *> O[2])=(0.0,0.0); 
        (A[6] *> O[3])=(0.0,0.0); 
        (A[6] *> O[4])=(0.0,0.0); 
        (A[6] *> O[5])=(0.0,0.0); 
        (A[6] *> O[6])=(0.0,0.0); 
        (A[6] *> O[7])=(0.0,0.0); 
        (A[6] *> O[8])=(0.0,0.0); 
        (A[6] *> O[9])=(0.0,0.0); 
        (A[6] *> O[10])=(0.0,0.0); 
        (A[6] *> O[11])=(0.0,0.0); 
        (A[6] *> O[12])=(0.0,0.0); 
        (A[6] *> O[13])=(0.0,0.0); 
        (A[6] *> O[14])=(0.0,0.0); 
        (A[6] *> O[15])=(0.0,0.0); 
        (A[6] *> O[16])=(0.0,0.0); 
        (A[6] *> O[17])=(0.0,0.0); 
        (A[6] *> O[18])=(0.0,0.0); 
        (A[6] *> O[19])=(0.0,0.0); 
        (A[6] *> O[20])=(0.0,0.0); 
        (A[6] *> O[21])=(0.0,0.0); 
        (A[6] *> O[22])=(0.0,0.0); 
        (A[6] *> O[23])=(0.0,0.0); 
        (A[6] *> O[24])=(0.0,0.0); 
        (A[6] *> O[25])=(0.0,0.0); 
        (A[6] *> O[26])=(0.0,0.0); 
        (A[6] *> O[27])=(0.0,0.0); 
        (A[6] *> O[28])=(0.0,0.0); 
        (A[6] *> O[29])=(0.0,0.0); 
        (A[6] *> O[30])=(0.0,0.0); 
        (A[6] *> O[31])=(0.0,0.0); 
        (A[7] *> O[0])=(0.0,0.0); 
        (A[7] *> O[1])=(0.0,0.0); 
        (A[7] *> O[2])=(0.0,0.0); 
        (A[7] *> O[3])=(0.0,0.0); 
        (A[7] *> O[4])=(0.0,0.0); 
        (A[7] *> O[5])=(0.0,0.0); 
        (A[7] *> O[6])=(0.0,0.0); 
        (A[7] *> O[7])=(0.0,0.0); 
        (A[7] *> O[8])=(0.0,0.0); 
        (A[7] *> O[9])=(0.0,0.0); 
        (A[7] *> O[10])=(0.0,0.0); 
        (A[7] *> O[11])=(0.0,0.0); 
        (A[7] *> O[12])=(0.0,0.0); 
        (A[7] *> O[13])=(0.0,0.0); 
        (A[7] *> O[14])=(0.0,0.0); 
        (A[7] *> O[15])=(0.0,0.0); 
        (A[7] *> O[16])=(0.0,0.0); 
        (A[7] *> O[17])=(0.0,0.0); 
        (A[7] *> O[18])=(0.0,0.0); 
        (A[7] *> O[19])=(0.0,0.0); 
        (A[7] *> O[20])=(0.0,0.0); 
        (A[7] *> O[21])=(0.0,0.0); 
        (A[7] *> O[22])=(0.0,0.0); 
        (A[7] *> O[23])=(0.0,0.0); 
        (A[7] *> O[24])=(0.0,0.0); 
        (A[7] *> O[25])=(0.0,0.0); 
        (A[7] *> O[26])=(0.0,0.0); 
        (A[7] *> O[27])=(0.0,0.0); 
        (A[7] *> O[28])=(0.0,0.0); 
        (A[7] *> O[29])=(0.0,0.0); 
        (A[7] *> O[30])=(0.0,0.0); 
        (A[7] *> O[31])=(0.0,0.0); 
        (A[8] *> O[0])=(0.0,0.0); 
        (A[8] *> O[1])=(0.0,0.0); 
        (A[8] *> O[2])=(0.0,0.0); 
        (A[8] *> O[3])=(0.0,0.0); 
        (A[8] *> O[4])=(0.0,0.0); 
        (A[8] *> O[5])=(0.0,0.0); 
        (A[8] *> O[6])=(0.0,0.0); 
        (A[8] *> O[7])=(0.0,0.0); 
        (A[8] *> O[8])=(0.0,0.0); 
        (A[8] *> O[9])=(0.0,0.0); 
        (A[8] *> O[10])=(0.0,0.0); 
        (A[8] *> O[11])=(0.0,0.0); 
        (A[8] *> O[12])=(0.0,0.0); 
        (A[8] *> O[13])=(0.0,0.0); 
        (A[8] *> O[14])=(0.0,0.0); 
        (A[8] *> O[15])=(0.0,0.0); 
        (A[8] *> O[16])=(0.0,0.0); 
        (A[8] *> O[17])=(0.0,0.0); 
        (A[8] *> O[18])=(0.0,0.0); 
        (A[8] *> O[19])=(0.0,0.0); 
        (A[8] *> O[20])=(0.0,0.0); 
        (A[8] *> O[21])=(0.0,0.0); 
        (A[8] *> O[22])=(0.0,0.0); 
        (A[8] *> O[23])=(0.0,0.0); 
        (A[8] *> O[24])=(0.0,0.0); 
        (A[8] *> O[25])=(0.0,0.0); 
        (A[8] *> O[26])=(0.0,0.0); 
        (A[8] *> O[27])=(0.0,0.0); 
        (A[8] *> O[28])=(0.0,0.0); 
        (A[8] *> O[29])=(0.0,0.0); 
        (A[8] *> O[30])=(0.0,0.0); 
        (A[8] *> O[31])=(0.0,0.0); 
        (A[9] *> O[0])=(0.0,0.0); 
        (A[9] *> O[1])=(0.0,0.0); 
        (A[9] *> O[2])=(0.0,0.0); 
        (A[9] *> O[3])=(0.0,0.0); 
        (A[9] *> O[4])=(0.0,0.0); 
        (A[9] *> O[5])=(0.0,0.0); 
        (A[9] *> O[6])=(0.0,0.0); 
        (A[9] *> O[7])=(0.0,0.0); 
        (A[9] *> O[8])=(0.0,0.0); 
        (A[9] *> O[9])=(0.0,0.0); 
        (A[9] *> O[10])=(0.0,0.0); 
        (A[9] *> O[11])=(0.0,0.0); 
        (A[9] *> O[12])=(0.0,0.0); 
        (A[9] *> O[13])=(0.0,0.0); 
        (A[9] *> O[14])=(0.0,0.0); 
        (A[9] *> O[15])=(0.0,0.0); 
        (A[9] *> O[16])=(0.0,0.0); 
        (A[9] *> O[17])=(0.0,0.0); 
        (A[9] *> O[18])=(0.0,0.0); 
        (A[9] *> O[19])=(0.0,0.0); 
        (A[9] *> O[20])=(0.0,0.0); 
        (A[9] *> O[21])=(0.0,0.0); 
        (A[9] *> O[22])=(0.0,0.0); 
        (A[9] *> O[23])=(0.0,0.0); 
        (A[9] *> O[24])=(0.0,0.0); 
        (A[9] *> O[25])=(0.0,0.0); 
        (A[9] *> O[26])=(0.0,0.0); 
        (A[9] *> O[27])=(0.0,0.0); 
        (A[9] *> O[28])=(0.0,0.0); 
        (A[9] *> O[29])=(0.0,0.0); 
        (A[9] *> O[30])=(0.0,0.0); 
        (A[9] *> O[31])=(0.0,0.0); 
        (A[10] *> O[0])=(0.0,0.0); 
        (A[10] *> O[1])=(0.0,0.0); 
        (A[10] *> O[2])=(0.0,0.0); 
        (A[10] *> O[3])=(0.0,0.0); 
        (A[10] *> O[4])=(0.0,0.0); 
        (A[10] *> O[5])=(0.0,0.0); 
        (A[10] *> O[6])=(0.0,0.0); 
        (A[10] *> O[7])=(0.0,0.0); 
        (A[10] *> O[8])=(0.0,0.0); 
        (A[10] *> O[9])=(0.0,0.0); 
        (A[10] *> O[10])=(0.0,0.0); 
        (A[10] *> O[11])=(0.0,0.0); 
        (A[10] *> O[12])=(0.0,0.0); 
        (A[10] *> O[13])=(0.0,0.0); 
        (A[10] *> O[14])=(0.0,0.0); 
        (A[10] *> O[15])=(0.0,0.0); 
        (A[10] *> O[16])=(0.0,0.0); 
        (A[10] *> O[17])=(0.0,0.0); 
        (A[10] *> O[18])=(0.0,0.0); 
        (A[10] *> O[19])=(0.0,0.0); 
        (A[10] *> O[20])=(0.0,0.0); 
        (A[10] *> O[21])=(0.0,0.0); 
        (A[10] *> O[22])=(0.0,0.0); 
        (A[10] *> O[23])=(0.0,0.0); 
        (A[10] *> O[24])=(0.0,0.0); 
        (A[10] *> O[25])=(0.0,0.0); 
        (A[10] *> O[26])=(0.0,0.0); 
        (A[10] *> O[27])=(0.0,0.0); 
        (A[10] *> O[28])=(0.0,0.0); 
        (A[10] *> O[29])=(0.0,0.0); 
        (A[10] *> O[30])=(0.0,0.0); 
        (A[10] *> O[31])=(0.0,0.0); 
        (A[11] *> O[0])=(0.0,0.0); 
        (A[11] *> O[1])=(0.0,0.0); 
        (A[11] *> O[2])=(0.0,0.0); 
        (A[11] *> O[3])=(0.0,0.0); 
        (A[11] *> O[4])=(0.0,0.0); 
        (A[11] *> O[5])=(0.0,0.0); 
        (A[11] *> O[6])=(0.0,0.0); 
        (A[11] *> O[7])=(0.0,0.0); 
        (A[11] *> O[8])=(0.0,0.0); 
        (A[11] *> O[9])=(0.0,0.0); 
        (A[11] *> O[10])=(0.0,0.0); 
        (A[11] *> O[11])=(0.0,0.0); 
        (A[11] *> O[12])=(0.0,0.0); 
        (A[11] *> O[13])=(0.0,0.0); 
        (A[11] *> O[14])=(0.0,0.0); 
        (A[11] *> O[15])=(0.0,0.0); 
        (A[11] *> O[16])=(0.0,0.0); 
        (A[11] *> O[17])=(0.0,0.0); 
        (A[11] *> O[18])=(0.0,0.0); 
        (A[11] *> O[19])=(0.0,0.0); 
        (A[11] *> O[20])=(0.0,0.0); 
        (A[11] *> O[21])=(0.0,0.0); 
        (A[11] *> O[22])=(0.0,0.0); 
        (A[11] *> O[23])=(0.0,0.0); 
        (A[11] *> O[24])=(0.0,0.0); 
        (A[11] *> O[25])=(0.0,0.0); 
        (A[11] *> O[26])=(0.0,0.0); 
        (A[11] *> O[27])=(0.0,0.0); 
        (A[11] *> O[28])=(0.0,0.0); 
        (A[11] *> O[29])=(0.0,0.0); 
        (A[11] *> O[30])=(0.0,0.0); 
        (A[11] *> O[31])=(0.0,0.0); 
        (A[12] *> O[0])=(0.0,0.0); 
        (A[12] *> O[1])=(0.0,0.0); 
        (A[12] *> O[2])=(0.0,0.0); 
        (A[12] *> O[3])=(0.0,0.0); 
        (A[12] *> O[4])=(0.0,0.0); 
        (A[12] *> O[5])=(0.0,0.0); 
        (A[12] *> O[6])=(0.0,0.0); 
        (A[12] *> O[7])=(0.0,0.0); 
        (A[12] *> O[8])=(0.0,0.0); 
        (A[12] *> O[9])=(0.0,0.0); 
        (A[12] *> O[10])=(0.0,0.0); 
        (A[12] *> O[11])=(0.0,0.0); 
        (A[12] *> O[12])=(0.0,0.0); 
        (A[12] *> O[13])=(0.0,0.0); 
        (A[12] *> O[14])=(0.0,0.0); 
        (A[12] *> O[15])=(0.0,0.0); 
        (A[12] *> O[16])=(0.0,0.0); 
        (A[12] *> O[17])=(0.0,0.0); 
        (A[12] *> O[18])=(0.0,0.0); 
        (A[12] *> O[19])=(0.0,0.0); 
        (A[12] *> O[20])=(0.0,0.0); 
        (A[12] *> O[21])=(0.0,0.0); 
        (A[12] *> O[22])=(0.0,0.0); 
        (A[12] *> O[23])=(0.0,0.0); 
        (A[12] *> O[24])=(0.0,0.0); 
        (A[12] *> O[25])=(0.0,0.0); 
        (A[12] *> O[26])=(0.0,0.0); 
        (A[12] *> O[27])=(0.0,0.0); 
        (A[12] *> O[28])=(0.0,0.0); 
        (A[12] *> O[29])=(0.0,0.0); 
        (A[12] *> O[30])=(0.0,0.0); 
        (A[12] *> O[31])=(0.0,0.0); 
        (A[13] *> O[0])=(0.0,0.0); 
        (A[13] *> O[1])=(0.0,0.0); 
        (A[13] *> O[2])=(0.0,0.0); 
        (A[13] *> O[3])=(0.0,0.0); 
        (A[13] *> O[4])=(0.0,0.0); 
        (A[13] *> O[5])=(0.0,0.0); 
        (A[13] *> O[6])=(0.0,0.0); 
        (A[13] *> O[7])=(0.0,0.0); 
        (A[13] *> O[8])=(0.0,0.0); 
        (A[13] *> O[9])=(0.0,0.0); 
        (A[13] *> O[10])=(0.0,0.0); 
        (A[13] *> O[11])=(0.0,0.0); 
        (A[13] *> O[12])=(0.0,0.0); 
        (A[13] *> O[13])=(0.0,0.0); 
        (A[13] *> O[14])=(0.0,0.0); 
        (A[13] *> O[15])=(0.0,0.0); 
        (A[13] *> O[16])=(0.0,0.0); 
        (A[13] *> O[17])=(0.0,0.0); 
        (A[13] *> O[18])=(0.0,0.0); 
        (A[13] *> O[19])=(0.0,0.0); 
        (A[13] *> O[20])=(0.0,0.0); 
        (A[13] *> O[21])=(0.0,0.0); 
        (A[13] *> O[22])=(0.0,0.0); 
        (A[13] *> O[23])=(0.0,0.0); 
        (A[13] *> O[24])=(0.0,0.0); 
        (A[13] *> O[25])=(0.0,0.0); 
        (A[13] *> O[26])=(0.0,0.0); 
        (A[13] *> O[27])=(0.0,0.0); 
        (A[13] *> O[28])=(0.0,0.0); 
        (A[13] *> O[29])=(0.0,0.0); 
        (A[13] *> O[30])=(0.0,0.0); 
        (A[13] *> O[31])=(0.0,0.0); 
        (A[14] *> O[0])=(0.0,0.0); 
        (A[14] *> O[1])=(0.0,0.0); 
        (A[14] *> O[2])=(0.0,0.0); 
        (A[14] *> O[3])=(0.0,0.0); 
        (A[14] *> O[4])=(0.0,0.0); 
        (A[14] *> O[5])=(0.0,0.0); 
        (A[14] *> O[6])=(0.0,0.0); 
        (A[14] *> O[7])=(0.0,0.0); 
        (A[14] *> O[8])=(0.0,0.0); 
        (A[14] *> O[9])=(0.0,0.0); 
        (A[14] *> O[10])=(0.0,0.0); 
        (A[14] *> O[11])=(0.0,0.0); 
        (A[14] *> O[12])=(0.0,0.0); 
        (A[14] *> O[13])=(0.0,0.0); 
        (A[14] *> O[14])=(0.0,0.0); 
        (A[14] *> O[15])=(0.0,0.0); 
        (A[14] *> O[16])=(0.0,0.0); 
        (A[14] *> O[17])=(0.0,0.0); 
        (A[14] *> O[18])=(0.0,0.0); 
        (A[14] *> O[19])=(0.0,0.0); 
        (A[14] *> O[20])=(0.0,0.0); 
        (A[14] *> O[21])=(0.0,0.0); 
        (A[14] *> O[22])=(0.0,0.0); 
        (A[14] *> O[23])=(0.0,0.0); 
        (A[14] *> O[24])=(0.0,0.0); 
        (A[14] *> O[25])=(0.0,0.0); 
        (A[14] *> O[26])=(0.0,0.0); 
        (A[14] *> O[27])=(0.0,0.0); 
        (A[14] *> O[28])=(0.0,0.0); 
        (A[14] *> O[29])=(0.0,0.0); 
        (A[14] *> O[30])=(0.0,0.0); 
        (A[14] *> O[31])=(0.0,0.0); 
        (A[15] *> O[0])=(0.0,0.0); 
        (A[15] *> O[1])=(0.0,0.0); 
        (A[15] *> O[2])=(0.0,0.0); 
        (A[15] *> O[3])=(0.0,0.0); 
        (A[15] *> O[4])=(0.0,0.0); 
        (A[15] *> O[5])=(0.0,0.0); 
        (A[15] *> O[6])=(0.0,0.0); 
        (A[15] *> O[7])=(0.0,0.0); 
        (A[15] *> O[8])=(0.0,0.0); 
        (A[15] *> O[9])=(0.0,0.0); 
        (A[15] *> O[10])=(0.0,0.0); 
        (A[15] *> O[11])=(0.0,0.0); 
        (A[15] *> O[12])=(0.0,0.0); 
        (A[15] *> O[13])=(0.0,0.0); 
        (A[15] *> O[14])=(0.0,0.0); 
        (A[15] *> O[15])=(0.0,0.0); 
        (A[15] *> O[16])=(0.0,0.0); 
        (A[15] *> O[17])=(0.0,0.0); 
        (A[15] *> O[18])=(0.0,0.0); 
        (A[15] *> O[19])=(0.0,0.0); 
        (A[15] *> O[20])=(0.0,0.0); 
        (A[15] *> O[21])=(0.0,0.0); 
        (A[15] *> O[22])=(0.0,0.0); 
        (A[15] *> O[23])=(0.0,0.0); 
        (A[15] *> O[24])=(0.0,0.0); 
        (A[15] *> O[25])=(0.0,0.0); 
        (A[15] *> O[26])=(0.0,0.0); 
        (A[15] *> O[27])=(0.0,0.0); 
        (A[15] *> O[28])=(0.0,0.0); 
        (A[15] *> O[29])=(0.0,0.0); 
        (A[15] *> O[30])=(0.0,0.0); 
        (A[15] *> O[31])=(0.0,0.0); 
        (B[0] *> O[0])=(0.0,0.0); 
        (B[0] *> O[1])=(0.0,0.0); 
        (B[0] *> O[2])=(0.0,0.0); 
        (B[0] *> O[3])=(0.0,0.0); 
        (B[0] *> O[4])=(0.0,0.0); 
        (B[0] *> O[5])=(0.0,0.0); 
        (B[0] *> O[6])=(0.0,0.0); 
        (B[0] *> O[7])=(0.0,0.0); 
        (B[0] *> O[8])=(0.0,0.0); 
        (B[0] *> O[9])=(0.0,0.0); 
        (B[0] *> O[10])=(0.0,0.0); 
        (B[0] *> O[11])=(0.0,0.0); 
        (B[0] *> O[12])=(0.0,0.0); 
        (B[0] *> O[13])=(0.0,0.0); 
        (B[0] *> O[14])=(0.0,0.0); 
        (B[0] *> O[15])=(0.0,0.0); 
        (B[0] *> O[16])=(0.0,0.0); 
        (B[0] *> O[17])=(0.0,0.0); 
        (B[0] *> O[18])=(0.0,0.0); 
        (B[0] *> O[19])=(0.0,0.0); 
        (B[0] *> O[20])=(0.0,0.0); 
        (B[0] *> O[21])=(0.0,0.0); 
        (B[0] *> O[22])=(0.0,0.0); 
        (B[0] *> O[23])=(0.0,0.0); 
        (B[0] *> O[24])=(0.0,0.0); 
        (B[0] *> O[25])=(0.0,0.0); 
        (B[0] *> O[26])=(0.0,0.0); 
        (B[0] *> O[27])=(0.0,0.0); 
        (B[0] *> O[28])=(0.0,0.0); 
        (B[0] *> O[29])=(0.0,0.0); 
        (B[0] *> O[30])=(0.0,0.0); 
        (B[0] *> O[31])=(0.0,0.0); 
        (B[1] *> O[0])=(0.0,0.0); 
        (B[1] *> O[1])=(0.0,0.0); 
        (B[1] *> O[2])=(0.0,0.0); 
        (B[1] *> O[3])=(0.0,0.0); 
        (B[1] *> O[4])=(0.0,0.0); 
        (B[1] *> O[5])=(0.0,0.0); 
        (B[1] *> O[6])=(0.0,0.0); 
        (B[1] *> O[7])=(0.0,0.0); 
        (B[1] *> O[8])=(0.0,0.0); 
        (B[1] *> O[9])=(0.0,0.0); 
        (B[1] *> O[10])=(0.0,0.0); 
        (B[1] *> O[11])=(0.0,0.0); 
        (B[1] *> O[12])=(0.0,0.0); 
        (B[1] *> O[13])=(0.0,0.0); 
        (B[1] *> O[14])=(0.0,0.0); 
        (B[1] *> O[15])=(0.0,0.0); 
        (B[1] *> O[16])=(0.0,0.0); 
        (B[1] *> O[17])=(0.0,0.0); 
        (B[1] *> O[18])=(0.0,0.0); 
        (B[1] *> O[19])=(0.0,0.0); 
        (B[1] *> O[20])=(0.0,0.0); 
        (B[1] *> O[21])=(0.0,0.0); 
        (B[1] *> O[22])=(0.0,0.0); 
        (B[1] *> O[23])=(0.0,0.0); 
        (B[1] *> O[24])=(0.0,0.0); 
        (B[1] *> O[25])=(0.0,0.0); 
        (B[1] *> O[26])=(0.0,0.0); 
        (B[1] *> O[27])=(0.0,0.0); 
        (B[1] *> O[28])=(0.0,0.0); 
        (B[1] *> O[29])=(0.0,0.0); 
        (B[1] *> O[30])=(0.0,0.0); 
        (B[1] *> O[31])=(0.0,0.0); 
        (B[2] *> O[0])=(0.0,0.0); 
        (B[2] *> O[1])=(0.0,0.0); 
        (B[2] *> O[2])=(0.0,0.0); 
        (B[2] *> O[3])=(0.0,0.0); 
        (B[2] *> O[4])=(0.0,0.0); 
        (B[2] *> O[5])=(0.0,0.0); 
        (B[2] *> O[6])=(0.0,0.0); 
        (B[2] *> O[7])=(0.0,0.0); 
        (B[2] *> O[8])=(0.0,0.0); 
        (B[2] *> O[9])=(0.0,0.0); 
        (B[2] *> O[10])=(0.0,0.0); 
        (B[2] *> O[11])=(0.0,0.0); 
        (B[2] *> O[12])=(0.0,0.0); 
        (B[2] *> O[13])=(0.0,0.0); 
        (B[2] *> O[14])=(0.0,0.0); 
        (B[2] *> O[15])=(0.0,0.0); 
        (B[2] *> O[16])=(0.0,0.0); 
        (B[2] *> O[17])=(0.0,0.0); 
        (B[2] *> O[18])=(0.0,0.0); 
        (B[2] *> O[19])=(0.0,0.0); 
        (B[2] *> O[20])=(0.0,0.0); 
        (B[2] *> O[21])=(0.0,0.0); 
        (B[2] *> O[22])=(0.0,0.0); 
        (B[2] *> O[23])=(0.0,0.0); 
        (B[2] *> O[24])=(0.0,0.0); 
        (B[2] *> O[25])=(0.0,0.0); 
        (B[2] *> O[26])=(0.0,0.0); 
        (B[2] *> O[27])=(0.0,0.0); 
        (B[2] *> O[28])=(0.0,0.0); 
        (B[2] *> O[29])=(0.0,0.0); 
        (B[2] *> O[30])=(0.0,0.0); 
        (B[2] *> O[31])=(0.0,0.0); 
        (B[3] *> O[0])=(0.0,0.0); 
        (B[3] *> O[1])=(0.0,0.0); 
        (B[3] *> O[2])=(0.0,0.0); 
        (B[3] *> O[3])=(0.0,0.0); 
        (B[3] *> O[4])=(0.0,0.0); 
        (B[3] *> O[5])=(0.0,0.0); 
        (B[3] *> O[6])=(0.0,0.0); 
        (B[3] *> O[7])=(0.0,0.0); 
        (B[3] *> O[8])=(0.0,0.0); 
        (B[3] *> O[9])=(0.0,0.0); 
        (B[3] *> O[10])=(0.0,0.0); 
        (B[3] *> O[11])=(0.0,0.0); 
        (B[3] *> O[12])=(0.0,0.0); 
        (B[3] *> O[13])=(0.0,0.0); 
        (B[3] *> O[14])=(0.0,0.0); 
        (B[3] *> O[15])=(0.0,0.0); 
        (B[3] *> O[16])=(0.0,0.0); 
        (B[3] *> O[17])=(0.0,0.0); 
        (B[3] *> O[18])=(0.0,0.0); 
        (B[3] *> O[19])=(0.0,0.0); 
        (B[3] *> O[20])=(0.0,0.0); 
        (B[3] *> O[21])=(0.0,0.0); 
        (B[3] *> O[22])=(0.0,0.0); 
        (B[3] *> O[23])=(0.0,0.0); 
        (B[3] *> O[24])=(0.0,0.0); 
        (B[3] *> O[25])=(0.0,0.0); 
        (B[3] *> O[26])=(0.0,0.0); 
        (B[3] *> O[27])=(0.0,0.0); 
        (B[3] *> O[28])=(0.0,0.0); 
        (B[3] *> O[29])=(0.0,0.0); 
        (B[3] *> O[30])=(0.0,0.0); 
        (B[3] *> O[31])=(0.0,0.0); 
        (B[4] *> O[0])=(0.0,0.0); 
        (B[4] *> O[1])=(0.0,0.0); 
        (B[4] *> O[2])=(0.0,0.0); 
        (B[4] *> O[3])=(0.0,0.0); 
        (B[4] *> O[4])=(0.0,0.0); 
        (B[4] *> O[5])=(0.0,0.0); 
        (B[4] *> O[6])=(0.0,0.0); 
        (B[4] *> O[7])=(0.0,0.0); 
        (B[4] *> O[8])=(0.0,0.0); 
        (B[4] *> O[9])=(0.0,0.0); 
        (B[4] *> O[10])=(0.0,0.0); 
        (B[4] *> O[11])=(0.0,0.0); 
        (B[4] *> O[12])=(0.0,0.0); 
        (B[4] *> O[13])=(0.0,0.0); 
        (B[4] *> O[14])=(0.0,0.0); 
        (B[4] *> O[15])=(0.0,0.0); 
        (B[4] *> O[16])=(0.0,0.0); 
        (B[4] *> O[17])=(0.0,0.0); 
        (B[4] *> O[18])=(0.0,0.0); 
        (B[4] *> O[19])=(0.0,0.0); 
        (B[4] *> O[20])=(0.0,0.0); 
        (B[4] *> O[21])=(0.0,0.0); 
        (B[4] *> O[22])=(0.0,0.0); 
        (B[4] *> O[23])=(0.0,0.0); 
        (B[4] *> O[24])=(0.0,0.0); 
        (B[4] *> O[25])=(0.0,0.0); 
        (B[4] *> O[26])=(0.0,0.0); 
        (B[4] *> O[27])=(0.0,0.0); 
        (B[4] *> O[28])=(0.0,0.0); 
        (B[4] *> O[29])=(0.0,0.0); 
        (B[4] *> O[30])=(0.0,0.0); 
        (B[4] *> O[31])=(0.0,0.0); 
        (B[5] *> O[0])=(0.0,0.0); 
        (B[5] *> O[1])=(0.0,0.0); 
        (B[5] *> O[2])=(0.0,0.0); 
        (B[5] *> O[3])=(0.0,0.0); 
        (B[5] *> O[4])=(0.0,0.0); 
        (B[5] *> O[5])=(0.0,0.0); 
        (B[5] *> O[6])=(0.0,0.0); 
        (B[5] *> O[7])=(0.0,0.0); 
        (B[5] *> O[8])=(0.0,0.0); 
        (B[5] *> O[9])=(0.0,0.0); 
        (B[5] *> O[10])=(0.0,0.0); 
        (B[5] *> O[11])=(0.0,0.0); 
        (B[5] *> O[12])=(0.0,0.0); 
        (B[5] *> O[13])=(0.0,0.0); 
        (B[5] *> O[14])=(0.0,0.0); 
        (B[5] *> O[15])=(0.0,0.0); 
        (B[5] *> O[16])=(0.0,0.0); 
        (B[5] *> O[17])=(0.0,0.0); 
        (B[5] *> O[18])=(0.0,0.0); 
        (B[5] *> O[19])=(0.0,0.0); 
        (B[5] *> O[20])=(0.0,0.0); 
        (B[5] *> O[21])=(0.0,0.0); 
        (B[5] *> O[22])=(0.0,0.0); 
        (B[5] *> O[23])=(0.0,0.0); 
        (B[5] *> O[24])=(0.0,0.0); 
        (B[5] *> O[25])=(0.0,0.0); 
        (B[5] *> O[26])=(0.0,0.0); 
        (B[5] *> O[27])=(0.0,0.0); 
        (B[5] *> O[28])=(0.0,0.0); 
        (B[5] *> O[29])=(0.0,0.0); 
        (B[5] *> O[30])=(0.0,0.0); 
        (B[5] *> O[31])=(0.0,0.0); 
        (B[6] *> O[0])=(0.0,0.0); 
        (B[6] *> O[1])=(0.0,0.0); 
        (B[6] *> O[2])=(0.0,0.0); 
        (B[6] *> O[3])=(0.0,0.0); 
        (B[6] *> O[4])=(0.0,0.0); 
        (B[6] *> O[5])=(0.0,0.0); 
        (B[6] *> O[6])=(0.0,0.0); 
        (B[6] *> O[7])=(0.0,0.0); 
        (B[6] *> O[8])=(0.0,0.0); 
        (B[6] *> O[9])=(0.0,0.0); 
        (B[6] *> O[10])=(0.0,0.0); 
        (B[6] *> O[11])=(0.0,0.0); 
        (B[6] *> O[12])=(0.0,0.0); 
        (B[6] *> O[13])=(0.0,0.0); 
        (B[6] *> O[14])=(0.0,0.0); 
        (B[6] *> O[15])=(0.0,0.0); 
        (B[6] *> O[16])=(0.0,0.0); 
        (B[6] *> O[17])=(0.0,0.0); 
        (B[6] *> O[18])=(0.0,0.0); 
        (B[6] *> O[19])=(0.0,0.0); 
        (B[6] *> O[20])=(0.0,0.0); 
        (B[6] *> O[21])=(0.0,0.0); 
        (B[6] *> O[22])=(0.0,0.0); 
        (B[6] *> O[23])=(0.0,0.0); 
        (B[6] *> O[24])=(0.0,0.0); 
        (B[6] *> O[25])=(0.0,0.0); 
        (B[6] *> O[26])=(0.0,0.0); 
        (B[6] *> O[27])=(0.0,0.0); 
        (B[6] *> O[28])=(0.0,0.0); 
        (B[6] *> O[29])=(0.0,0.0); 
        (B[6] *> O[30])=(0.0,0.0); 
        (B[6] *> O[31])=(0.0,0.0); 
        (B[7] *> O[0])=(0.0,0.0); 
        (B[7] *> O[1])=(0.0,0.0); 
        (B[7] *> O[2])=(0.0,0.0); 
        (B[7] *> O[3])=(0.0,0.0); 
        (B[7] *> O[4])=(0.0,0.0); 
        (B[7] *> O[5])=(0.0,0.0); 
        (B[7] *> O[6])=(0.0,0.0); 
        (B[7] *> O[7])=(0.0,0.0); 
        (B[7] *> O[8])=(0.0,0.0); 
        (B[7] *> O[9])=(0.0,0.0); 
        (B[7] *> O[10])=(0.0,0.0); 
        (B[7] *> O[11])=(0.0,0.0); 
        (B[7] *> O[12])=(0.0,0.0); 
        (B[7] *> O[13])=(0.0,0.0); 
        (B[7] *> O[14])=(0.0,0.0); 
        (B[7] *> O[15])=(0.0,0.0); 
        (B[7] *> O[16])=(0.0,0.0); 
        (B[7] *> O[17])=(0.0,0.0); 
        (B[7] *> O[18])=(0.0,0.0); 
        (B[7] *> O[19])=(0.0,0.0); 
        (B[7] *> O[20])=(0.0,0.0); 
        (B[7] *> O[21])=(0.0,0.0); 
        (B[7] *> O[22])=(0.0,0.0); 
        (B[7] *> O[23])=(0.0,0.0); 
        (B[7] *> O[24])=(0.0,0.0); 
        (B[7] *> O[25])=(0.0,0.0); 
        (B[7] *> O[26])=(0.0,0.0); 
        (B[7] *> O[27])=(0.0,0.0); 
        (B[7] *> O[28])=(0.0,0.0); 
        (B[7] *> O[29])=(0.0,0.0); 
        (B[7] *> O[30])=(0.0,0.0); 
        (B[7] *> O[31])=(0.0,0.0); 
        (B[8] *> O[0])=(0.0,0.0); 
        (B[8] *> O[1])=(0.0,0.0); 
        (B[8] *> O[2])=(0.0,0.0); 
        (B[8] *> O[3])=(0.0,0.0); 
        (B[8] *> O[4])=(0.0,0.0); 
        (B[8] *> O[5])=(0.0,0.0); 
        (B[8] *> O[6])=(0.0,0.0); 
        (B[8] *> O[7])=(0.0,0.0); 
        (B[8] *> O[8])=(0.0,0.0); 
        (B[8] *> O[9])=(0.0,0.0); 
        (B[8] *> O[10])=(0.0,0.0); 
        (B[8] *> O[11])=(0.0,0.0); 
        (B[8] *> O[12])=(0.0,0.0); 
        (B[8] *> O[13])=(0.0,0.0); 
        (B[8] *> O[14])=(0.0,0.0); 
        (B[8] *> O[15])=(0.0,0.0); 
        (B[8] *> O[16])=(0.0,0.0); 
        (B[8] *> O[17])=(0.0,0.0); 
        (B[8] *> O[18])=(0.0,0.0); 
        (B[8] *> O[19])=(0.0,0.0); 
        (B[8] *> O[20])=(0.0,0.0); 
        (B[8] *> O[21])=(0.0,0.0); 
        (B[8] *> O[22])=(0.0,0.0); 
        (B[8] *> O[23])=(0.0,0.0); 
        (B[8] *> O[24])=(0.0,0.0); 
        (B[8] *> O[25])=(0.0,0.0); 
        (B[8] *> O[26])=(0.0,0.0); 
        (B[8] *> O[27])=(0.0,0.0); 
        (B[8] *> O[28])=(0.0,0.0); 
        (B[8] *> O[29])=(0.0,0.0); 
        (B[8] *> O[30])=(0.0,0.0); 
        (B[8] *> O[31])=(0.0,0.0); 
        (B[9] *> O[0])=(0.0,0.0); 
        (B[9] *> O[1])=(0.0,0.0); 
        (B[9] *> O[2])=(0.0,0.0); 
        (B[9] *> O[3])=(0.0,0.0); 
        (B[9] *> O[4])=(0.0,0.0); 
        (B[9] *> O[5])=(0.0,0.0); 
        (B[9] *> O[6])=(0.0,0.0); 
        (B[9] *> O[7])=(0.0,0.0); 
        (B[9] *> O[8])=(0.0,0.0); 
        (B[9] *> O[9])=(0.0,0.0); 
        (B[9] *> O[10])=(0.0,0.0); 
        (B[9] *> O[11])=(0.0,0.0); 
        (B[9] *> O[12])=(0.0,0.0); 
        (B[9] *> O[13])=(0.0,0.0); 
        (B[9] *> O[14])=(0.0,0.0); 
        (B[9] *> O[15])=(0.0,0.0); 
        (B[9] *> O[16])=(0.0,0.0); 
        (B[9] *> O[17])=(0.0,0.0); 
        (B[9] *> O[18])=(0.0,0.0); 
        (B[9] *> O[19])=(0.0,0.0); 
        (B[9] *> O[20])=(0.0,0.0); 
        (B[9] *> O[21])=(0.0,0.0); 
        (B[9] *> O[22])=(0.0,0.0); 
        (B[9] *> O[23])=(0.0,0.0); 
        (B[9] *> O[24])=(0.0,0.0); 
        (B[9] *> O[25])=(0.0,0.0); 
        (B[9] *> O[26])=(0.0,0.0); 
        (B[9] *> O[27])=(0.0,0.0); 
        (B[9] *> O[28])=(0.0,0.0); 
        (B[9] *> O[29])=(0.0,0.0); 
        (B[9] *> O[30])=(0.0,0.0); 
        (B[9] *> O[31])=(0.0,0.0); 
        (B[10] *> O[0])=(0.0,0.0); 
        (B[10] *> O[1])=(0.0,0.0); 
        (B[10] *> O[2])=(0.0,0.0); 
        (B[10] *> O[3])=(0.0,0.0); 
        (B[10] *> O[4])=(0.0,0.0); 
        (B[10] *> O[5])=(0.0,0.0); 
        (B[10] *> O[6])=(0.0,0.0); 
        (B[10] *> O[7])=(0.0,0.0); 
        (B[10] *> O[8])=(0.0,0.0); 
        (B[10] *> O[9])=(0.0,0.0); 
        (B[10] *> O[10])=(0.0,0.0); 
        (B[10] *> O[11])=(0.0,0.0); 
        (B[10] *> O[12])=(0.0,0.0); 
        (B[10] *> O[13])=(0.0,0.0); 
        (B[10] *> O[14])=(0.0,0.0); 
        (B[10] *> O[15])=(0.0,0.0); 
        (B[10] *> O[16])=(0.0,0.0); 
        (B[10] *> O[17])=(0.0,0.0); 
        (B[10] *> O[18])=(0.0,0.0); 
        (B[10] *> O[19])=(0.0,0.0); 
        (B[10] *> O[20])=(0.0,0.0); 
        (B[10] *> O[21])=(0.0,0.0); 
        (B[10] *> O[22])=(0.0,0.0); 
        (B[10] *> O[23])=(0.0,0.0); 
        (B[10] *> O[24])=(0.0,0.0); 
        (B[10] *> O[25])=(0.0,0.0); 
        (B[10] *> O[26])=(0.0,0.0); 
        (B[10] *> O[27])=(0.0,0.0); 
        (B[10] *> O[28])=(0.0,0.0); 
        (B[10] *> O[29])=(0.0,0.0); 
        (B[10] *> O[30])=(0.0,0.0); 
        (B[10] *> O[31])=(0.0,0.0); 
        (B[11] *> O[0])=(0.0,0.0); 
        (B[11] *> O[1])=(0.0,0.0); 
        (B[11] *> O[2])=(0.0,0.0); 
        (B[11] *> O[3])=(0.0,0.0); 
        (B[11] *> O[4])=(0.0,0.0); 
        (B[11] *> O[5])=(0.0,0.0); 
        (B[11] *> O[6])=(0.0,0.0); 
        (B[11] *> O[7])=(0.0,0.0); 
        (B[11] *> O[8])=(0.0,0.0); 
        (B[11] *> O[9])=(0.0,0.0); 
        (B[11] *> O[10])=(0.0,0.0); 
        (B[11] *> O[11])=(0.0,0.0); 
        (B[11] *> O[12])=(0.0,0.0); 
        (B[11] *> O[13])=(0.0,0.0); 
        (B[11] *> O[14])=(0.0,0.0); 
        (B[11] *> O[15])=(0.0,0.0); 
        (B[11] *> O[16])=(0.0,0.0); 
        (B[11] *> O[17])=(0.0,0.0); 
        (B[11] *> O[18])=(0.0,0.0); 
        (B[11] *> O[19])=(0.0,0.0); 
        (B[11] *> O[20])=(0.0,0.0); 
        (B[11] *> O[21])=(0.0,0.0); 
        (B[11] *> O[22])=(0.0,0.0); 
        (B[11] *> O[23])=(0.0,0.0); 
        (B[11] *> O[24])=(0.0,0.0); 
        (B[11] *> O[25])=(0.0,0.0); 
        (B[11] *> O[26])=(0.0,0.0); 
        (B[11] *> O[27])=(0.0,0.0); 
        (B[11] *> O[28])=(0.0,0.0); 
        (B[11] *> O[29])=(0.0,0.0); 
        (B[11] *> O[30])=(0.0,0.0); 
        (B[11] *> O[31])=(0.0,0.0); 
        (B[12] *> O[0])=(0.0,0.0); 
        (B[12] *> O[1])=(0.0,0.0); 
        (B[12] *> O[2])=(0.0,0.0); 
        (B[12] *> O[3])=(0.0,0.0); 
        (B[12] *> O[4])=(0.0,0.0); 
        (B[12] *> O[5])=(0.0,0.0); 
        (B[12] *> O[6])=(0.0,0.0); 
        (B[12] *> O[7])=(0.0,0.0); 
        (B[12] *> O[8])=(0.0,0.0); 
        (B[12] *> O[9])=(0.0,0.0); 
        (B[12] *> O[10])=(0.0,0.0); 
        (B[12] *> O[11])=(0.0,0.0); 
        (B[12] *> O[12])=(0.0,0.0); 
        (B[12] *> O[13])=(0.0,0.0); 
        (B[12] *> O[14])=(0.0,0.0); 
        (B[12] *> O[15])=(0.0,0.0); 
        (B[12] *> O[16])=(0.0,0.0); 
        (B[12] *> O[17])=(0.0,0.0); 
        (B[12] *> O[18])=(0.0,0.0); 
        (B[12] *> O[19])=(0.0,0.0); 
        (B[12] *> O[20])=(0.0,0.0); 
        (B[12] *> O[21])=(0.0,0.0); 
        (B[12] *> O[22])=(0.0,0.0); 
        (B[12] *> O[23])=(0.0,0.0); 
        (B[12] *> O[24])=(0.0,0.0); 
        (B[12] *> O[25])=(0.0,0.0); 
        (B[12] *> O[26])=(0.0,0.0); 
        (B[12] *> O[27])=(0.0,0.0); 
        (B[12] *> O[28])=(0.0,0.0); 
        (B[12] *> O[29])=(0.0,0.0); 
        (B[12] *> O[30])=(0.0,0.0); 
        (B[12] *> O[31])=(0.0,0.0); 
        (B[13] *> O[0])=(0.0,0.0); 
        (B[13] *> O[1])=(0.0,0.0); 
        (B[13] *> O[2])=(0.0,0.0); 
        (B[13] *> O[3])=(0.0,0.0); 
        (B[13] *> O[4])=(0.0,0.0); 
        (B[13] *> O[5])=(0.0,0.0); 
        (B[13] *> O[6])=(0.0,0.0); 
        (B[13] *> O[7])=(0.0,0.0); 
        (B[13] *> O[8])=(0.0,0.0); 
        (B[13] *> O[9])=(0.0,0.0); 
        (B[13] *> O[10])=(0.0,0.0); 
        (B[13] *> O[11])=(0.0,0.0); 
        (B[13] *> O[12])=(0.0,0.0); 
        (B[13] *> O[13])=(0.0,0.0); 
        (B[13] *> O[14])=(0.0,0.0); 
        (B[13] *> O[15])=(0.0,0.0); 
        (B[13] *> O[16])=(0.0,0.0); 
        (B[13] *> O[17])=(0.0,0.0); 
        (B[13] *> O[18])=(0.0,0.0); 
        (B[13] *> O[19])=(0.0,0.0); 
        (B[13] *> O[20])=(0.0,0.0); 
        (B[13] *> O[21])=(0.0,0.0); 
        (B[13] *> O[22])=(0.0,0.0); 
        (B[13] *> O[23])=(0.0,0.0); 
        (B[13] *> O[24])=(0.0,0.0); 
        (B[13] *> O[25])=(0.0,0.0); 
        (B[13] *> O[26])=(0.0,0.0); 
        (B[13] *> O[27])=(0.0,0.0); 
        (B[13] *> O[28])=(0.0,0.0); 
        (B[13] *> O[29])=(0.0,0.0); 
        (B[13] *> O[30])=(0.0,0.0); 
        (B[13] *> O[31])=(0.0,0.0); 
        (B[14] *> O[0])=(0.0,0.0); 
        (B[14] *> O[1])=(0.0,0.0); 
        (B[14] *> O[2])=(0.0,0.0); 
        (B[14] *> O[3])=(0.0,0.0); 
        (B[14] *> O[4])=(0.0,0.0); 
        (B[14] *> O[5])=(0.0,0.0); 
        (B[14] *> O[6])=(0.0,0.0); 
        (B[14] *> O[7])=(0.0,0.0); 
        (B[14] *> O[8])=(0.0,0.0); 
        (B[14] *> O[9])=(0.0,0.0); 
        (B[14] *> O[10])=(0.0,0.0); 
        (B[14] *> O[11])=(0.0,0.0); 
        (B[14] *> O[12])=(0.0,0.0); 
        (B[14] *> O[13])=(0.0,0.0); 
        (B[14] *> O[14])=(0.0,0.0); 
        (B[14] *> O[15])=(0.0,0.0); 
        (B[14] *> O[16])=(0.0,0.0); 
        (B[14] *> O[17])=(0.0,0.0); 
        (B[14] *> O[18])=(0.0,0.0); 
        (B[14] *> O[19])=(0.0,0.0); 
        (B[14] *> O[20])=(0.0,0.0); 
        (B[14] *> O[21])=(0.0,0.0); 
        (B[14] *> O[22])=(0.0,0.0); 
        (B[14] *> O[23])=(0.0,0.0); 
        (B[14] *> O[24])=(0.0,0.0); 
        (B[14] *> O[25])=(0.0,0.0); 
        (B[14] *> O[26])=(0.0,0.0); 
        (B[14] *> O[27])=(0.0,0.0); 
        (B[14] *> O[28])=(0.0,0.0); 
        (B[14] *> O[29])=(0.0,0.0); 
        (B[14] *> O[30])=(0.0,0.0); 
        (B[14] *> O[31])=(0.0,0.0); 
        (B[15] *> O[0])=(0.0,0.0); 
        (B[15] *> O[1])=(0.0,0.0); 
        (B[15] *> O[2])=(0.0,0.0); 
        (B[15] *> O[3])=(0.0,0.0); 
        (B[15] *> O[4])=(0.0,0.0); 
        (B[15] *> O[5])=(0.0,0.0); 
        (B[15] *> O[6])=(0.0,0.0); 
        (B[15] *> O[7])=(0.0,0.0); 
        (B[15] *> O[8])=(0.0,0.0); 
        (B[15] *> O[9])=(0.0,0.0); 
        (B[15] *> O[10])=(0.0,0.0); 
        (B[15] *> O[11])=(0.0,0.0); 
        (B[15] *> O[12])=(0.0,0.0); 
        (B[15] *> O[13])=(0.0,0.0); 
        (B[15] *> O[14])=(0.0,0.0); 
        (B[15] *> O[15])=(0.0,0.0); 
        (B[15] *> O[16])=(0.0,0.0); 
        (B[15] *> O[17])=(0.0,0.0); 
        (B[15] *> O[18])=(0.0,0.0); 
        (B[15] *> O[19])=(0.0,0.0); 
        (B[15] *> O[20])=(0.0,0.0); 
        (B[15] *> O[21])=(0.0,0.0); 
        (B[15] *> O[22])=(0.0,0.0); 
        (B[15] *> O[23])=(0.0,0.0); 
        (B[15] *> O[24])=(0.0,0.0); 
        (B[15] *> O[25])=(0.0,0.0); 
        (B[15] *> O[26])=(0.0,0.0); 
        (B[15] *> O[27])=(0.0,0.0); 
        (B[15] *> O[28])=(0.0,0.0); 
        (B[15] *> O[29])=(0.0,0.0); 
        (B[15] *> O[30])=(0.0,0.0); 
        (B[15] *> O[31])=(0.0,0.0); 
        (C[0] *> O[0])=(0.0,0.0); 
        (C[0] *> O[1])=(0.0,0.0); 
        (C[0] *> O[2])=(0.0,0.0); 
        (C[0] *> O[3])=(0.0,0.0); 
        (C[0] *> O[4])=(0.0,0.0); 
        (C[0] *> O[5])=(0.0,0.0); 
        (C[0] *> O[6])=(0.0,0.0); 
        (C[0] *> O[7])=(0.0,0.0); 
        (C[0] *> O[8])=(0.0,0.0); 
        (C[0] *> O[9])=(0.0,0.0); 
        (C[0] *> O[10])=(0.0,0.0); 
        (C[0] *> O[11])=(0.0,0.0); 
        (C[0] *> O[12])=(0.0,0.0); 
        (C[0] *> O[13])=(0.0,0.0); 
        (C[0] *> O[14])=(0.0,0.0); 
        (C[0] *> O[15])=(0.0,0.0); 
        (C[0] *> O[16])=(0.0,0.0); 
        (C[0] *> O[17])=(0.0,0.0); 
        (C[0] *> O[18])=(0.0,0.0); 
        (C[0] *> O[19])=(0.0,0.0); 
        (C[0] *> O[20])=(0.0,0.0); 
        (C[0] *> O[21])=(0.0,0.0); 
        (C[0] *> O[22])=(0.0,0.0); 
        (C[0] *> O[23])=(0.0,0.0); 
        (C[0] *> O[24])=(0.0,0.0); 
        (C[0] *> O[25])=(0.0,0.0); 
        (C[0] *> O[26])=(0.0,0.0); 
        (C[0] *> O[27])=(0.0,0.0); 
        (C[0] *> O[28])=(0.0,0.0); 
        (C[0] *> O[29])=(0.0,0.0); 
        (C[0] *> O[30])=(0.0,0.0); 
        (C[0] *> O[31])=(0.0,0.0); 
        (C[1] *> O[0])=(0.0,0.0); 
        (C[1] *> O[1])=(0.0,0.0); 
        (C[1] *> O[2])=(0.0,0.0); 
        (C[1] *> O[3])=(0.0,0.0); 
        (C[1] *> O[4])=(0.0,0.0); 
        (C[1] *> O[5])=(0.0,0.0); 
        (C[1] *> O[6])=(0.0,0.0); 
        (C[1] *> O[7])=(0.0,0.0); 
        (C[1] *> O[8])=(0.0,0.0); 
        (C[1] *> O[9])=(0.0,0.0); 
        (C[1] *> O[10])=(0.0,0.0); 
        (C[1] *> O[11])=(0.0,0.0); 
        (C[1] *> O[12])=(0.0,0.0); 
        (C[1] *> O[13])=(0.0,0.0); 
        (C[1] *> O[14])=(0.0,0.0); 
        (C[1] *> O[15])=(0.0,0.0); 
        (C[1] *> O[16])=(0.0,0.0); 
        (C[1] *> O[17])=(0.0,0.0); 
        (C[1] *> O[18])=(0.0,0.0); 
        (C[1] *> O[19])=(0.0,0.0); 
        (C[1] *> O[20])=(0.0,0.0); 
        (C[1] *> O[21])=(0.0,0.0); 
        (C[1] *> O[22])=(0.0,0.0); 
        (C[1] *> O[23])=(0.0,0.0); 
        (C[1] *> O[24])=(0.0,0.0); 
        (C[1] *> O[25])=(0.0,0.0); 
        (C[1] *> O[26])=(0.0,0.0); 
        (C[1] *> O[27])=(0.0,0.0); 
        (C[1] *> O[28])=(0.0,0.0); 
        (C[1] *> O[29])=(0.0,0.0); 
        (C[1] *> O[30])=(0.0,0.0); 
        (C[1] *> O[31])=(0.0,0.0); 
        (C[2] *> O[0])=(0.0,0.0); 
        (C[2] *> O[1])=(0.0,0.0); 
        (C[2] *> O[2])=(0.0,0.0); 
        (C[2] *> O[3])=(0.0,0.0); 
        (C[2] *> O[4])=(0.0,0.0); 
        (C[2] *> O[5])=(0.0,0.0); 
        (C[2] *> O[6])=(0.0,0.0); 
        (C[2] *> O[7])=(0.0,0.0); 
        (C[2] *> O[8])=(0.0,0.0); 
        (C[2] *> O[9])=(0.0,0.0); 
        (C[2] *> O[10])=(0.0,0.0); 
        (C[2] *> O[11])=(0.0,0.0); 
        (C[2] *> O[12])=(0.0,0.0); 
        (C[2] *> O[13])=(0.0,0.0); 
        (C[2] *> O[14])=(0.0,0.0); 
        (C[2] *> O[15])=(0.0,0.0); 
        (C[2] *> O[16])=(0.0,0.0); 
        (C[2] *> O[17])=(0.0,0.0); 
        (C[2] *> O[18])=(0.0,0.0); 
        (C[2] *> O[19])=(0.0,0.0); 
        (C[2] *> O[20])=(0.0,0.0); 
        (C[2] *> O[21])=(0.0,0.0); 
        (C[2] *> O[22])=(0.0,0.0); 
        (C[2] *> O[23])=(0.0,0.0); 
        (C[2] *> O[24])=(0.0,0.0); 
        (C[2] *> O[25])=(0.0,0.0); 
        (C[2] *> O[26])=(0.0,0.0); 
        (C[2] *> O[27])=(0.0,0.0); 
        (C[2] *> O[28])=(0.0,0.0); 
        (C[2] *> O[29])=(0.0,0.0); 
        (C[2] *> O[30])=(0.0,0.0); 
        (C[2] *> O[31])=(0.0,0.0); 
        (C[3] *> O[0])=(0.0,0.0); 
        (C[3] *> O[1])=(0.0,0.0); 
        (C[3] *> O[2])=(0.0,0.0); 
        (C[3] *> O[3])=(0.0,0.0); 
        (C[3] *> O[4])=(0.0,0.0); 
        (C[3] *> O[5])=(0.0,0.0); 
        (C[3] *> O[6])=(0.0,0.0); 
        (C[3] *> O[7])=(0.0,0.0); 
        (C[3] *> O[8])=(0.0,0.0); 
        (C[3] *> O[9])=(0.0,0.0); 
        (C[3] *> O[10])=(0.0,0.0); 
        (C[3] *> O[11])=(0.0,0.0); 
        (C[3] *> O[12])=(0.0,0.0); 
        (C[3] *> O[13])=(0.0,0.0); 
        (C[3] *> O[14])=(0.0,0.0); 
        (C[3] *> O[15])=(0.0,0.0); 
        (C[3] *> O[16])=(0.0,0.0); 
        (C[3] *> O[17])=(0.0,0.0); 
        (C[3] *> O[18])=(0.0,0.0); 
        (C[3] *> O[19])=(0.0,0.0); 
        (C[3] *> O[20])=(0.0,0.0); 
        (C[3] *> O[21])=(0.0,0.0); 
        (C[3] *> O[22])=(0.0,0.0); 
        (C[3] *> O[23])=(0.0,0.0); 
        (C[3] *> O[24])=(0.0,0.0); 
        (C[3] *> O[25])=(0.0,0.0); 
        (C[3] *> O[26])=(0.0,0.0); 
        (C[3] *> O[27])=(0.0,0.0); 
        (C[3] *> O[28])=(0.0,0.0); 
        (C[3] *> O[29])=(0.0,0.0); 
        (C[3] *> O[30])=(0.0,0.0); 
        (C[3] *> O[31])=(0.0,0.0); 
        (C[4] *> O[0])=(0.0,0.0); 
        (C[4] *> O[1])=(0.0,0.0); 
        (C[4] *> O[2])=(0.0,0.0); 
        (C[4] *> O[3])=(0.0,0.0); 
        (C[4] *> O[4])=(0.0,0.0); 
        (C[4] *> O[5])=(0.0,0.0); 
        (C[4] *> O[6])=(0.0,0.0); 
        (C[4] *> O[7])=(0.0,0.0); 
        (C[4] *> O[8])=(0.0,0.0); 
        (C[4] *> O[9])=(0.0,0.0); 
        (C[4] *> O[10])=(0.0,0.0); 
        (C[4] *> O[11])=(0.0,0.0); 
        (C[4] *> O[12])=(0.0,0.0); 
        (C[4] *> O[13])=(0.0,0.0); 
        (C[4] *> O[14])=(0.0,0.0); 
        (C[4] *> O[15])=(0.0,0.0); 
        (C[4] *> O[16])=(0.0,0.0); 
        (C[4] *> O[17])=(0.0,0.0); 
        (C[4] *> O[18])=(0.0,0.0); 
        (C[4] *> O[19])=(0.0,0.0); 
        (C[4] *> O[20])=(0.0,0.0); 
        (C[4] *> O[21])=(0.0,0.0); 
        (C[4] *> O[22])=(0.0,0.0); 
        (C[4] *> O[23])=(0.0,0.0); 
        (C[4] *> O[24])=(0.0,0.0); 
        (C[4] *> O[25])=(0.0,0.0); 
        (C[4] *> O[26])=(0.0,0.0); 
        (C[4] *> O[27])=(0.0,0.0); 
        (C[4] *> O[28])=(0.0,0.0); 
        (C[4] *> O[29])=(0.0,0.0); 
        (C[4] *> O[30])=(0.0,0.0); 
        (C[4] *> O[31])=(0.0,0.0); 
        (C[5] *> O[0])=(0.0,0.0); 
        (C[5] *> O[1])=(0.0,0.0); 
        (C[5] *> O[2])=(0.0,0.0); 
        (C[5] *> O[3])=(0.0,0.0); 
        (C[5] *> O[4])=(0.0,0.0); 
        (C[5] *> O[5])=(0.0,0.0); 
        (C[5] *> O[6])=(0.0,0.0); 
        (C[5] *> O[7])=(0.0,0.0); 
        (C[5] *> O[8])=(0.0,0.0); 
        (C[5] *> O[9])=(0.0,0.0); 
        (C[5] *> O[10])=(0.0,0.0); 
        (C[5] *> O[11])=(0.0,0.0); 
        (C[5] *> O[12])=(0.0,0.0); 
        (C[5] *> O[13])=(0.0,0.0); 
        (C[5] *> O[14])=(0.0,0.0); 
        (C[5] *> O[15])=(0.0,0.0); 
        (C[5] *> O[16])=(0.0,0.0); 
        (C[5] *> O[17])=(0.0,0.0); 
        (C[5] *> O[18])=(0.0,0.0); 
        (C[5] *> O[19])=(0.0,0.0); 
        (C[5] *> O[20])=(0.0,0.0); 
        (C[5] *> O[21])=(0.0,0.0); 
        (C[5] *> O[22])=(0.0,0.0); 
        (C[5] *> O[23])=(0.0,0.0); 
        (C[5] *> O[24])=(0.0,0.0); 
        (C[5] *> O[25])=(0.0,0.0); 
        (C[5] *> O[26])=(0.0,0.0); 
        (C[5] *> O[27])=(0.0,0.0); 
        (C[5] *> O[28])=(0.0,0.0); 
        (C[5] *> O[29])=(0.0,0.0); 
        (C[5] *> O[30])=(0.0,0.0); 
        (C[5] *> O[31])=(0.0,0.0); 
        (C[6] *> O[0])=(0.0,0.0); 
        (C[6] *> O[1])=(0.0,0.0); 
        (C[6] *> O[2])=(0.0,0.0); 
        (C[6] *> O[3])=(0.0,0.0); 
        (C[6] *> O[4])=(0.0,0.0); 
        (C[6] *> O[5])=(0.0,0.0); 
        (C[6] *> O[6])=(0.0,0.0); 
        (C[6] *> O[7])=(0.0,0.0); 
        (C[6] *> O[8])=(0.0,0.0); 
        (C[6] *> O[9])=(0.0,0.0); 
        (C[6] *> O[10])=(0.0,0.0); 
        (C[6] *> O[11])=(0.0,0.0); 
        (C[6] *> O[12])=(0.0,0.0); 
        (C[6] *> O[13])=(0.0,0.0); 
        (C[6] *> O[14])=(0.0,0.0); 
        (C[6] *> O[15])=(0.0,0.0); 
        (C[6] *> O[16])=(0.0,0.0); 
        (C[6] *> O[17])=(0.0,0.0); 
        (C[6] *> O[18])=(0.0,0.0); 
        (C[6] *> O[19])=(0.0,0.0); 
        (C[6] *> O[20])=(0.0,0.0); 
        (C[6] *> O[21])=(0.0,0.0); 
        (C[6] *> O[22])=(0.0,0.0); 
        (C[6] *> O[23])=(0.0,0.0); 
        (C[6] *> O[24])=(0.0,0.0); 
        (C[6] *> O[25])=(0.0,0.0); 
        (C[6] *> O[26])=(0.0,0.0); 
        (C[6] *> O[27])=(0.0,0.0); 
        (C[6] *> O[28])=(0.0,0.0); 
        (C[6] *> O[29])=(0.0,0.0); 
        (C[6] *> O[30])=(0.0,0.0); 
        (C[6] *> O[31])=(0.0,0.0); 
        (C[7] *> O[0])=(0.0,0.0); 
        (C[7] *> O[1])=(0.0,0.0); 
        (C[7] *> O[2])=(0.0,0.0); 
        (C[7] *> O[3])=(0.0,0.0); 
        (C[7] *> O[4])=(0.0,0.0); 
        (C[7] *> O[5])=(0.0,0.0); 
        (C[7] *> O[6])=(0.0,0.0); 
        (C[7] *> O[7])=(0.0,0.0); 
        (C[7] *> O[8])=(0.0,0.0); 
        (C[7] *> O[9])=(0.0,0.0); 
        (C[7] *> O[10])=(0.0,0.0); 
        (C[7] *> O[11])=(0.0,0.0); 
        (C[7] *> O[12])=(0.0,0.0); 
        (C[7] *> O[13])=(0.0,0.0); 
        (C[7] *> O[14])=(0.0,0.0); 
        (C[7] *> O[15])=(0.0,0.0); 
        (C[7] *> O[16])=(0.0,0.0); 
        (C[7] *> O[17])=(0.0,0.0); 
        (C[7] *> O[18])=(0.0,0.0); 
        (C[7] *> O[19])=(0.0,0.0); 
        (C[7] *> O[20])=(0.0,0.0); 
        (C[7] *> O[21])=(0.0,0.0); 
        (C[7] *> O[22])=(0.0,0.0); 
        (C[7] *> O[23])=(0.0,0.0); 
        (C[7] *> O[24])=(0.0,0.0); 
        (C[7] *> O[25])=(0.0,0.0); 
        (C[7] *> O[26])=(0.0,0.0); 
        (C[7] *> O[27])=(0.0,0.0); 
        (C[7] *> O[28])=(0.0,0.0); 
        (C[7] *> O[29])=(0.0,0.0); 
        (C[7] *> O[30])=(0.0,0.0); 
        (C[7] *> O[31])=(0.0,0.0); 
        (C[8] *> O[0])=(0.0,0.0); 
        (C[8] *> O[1])=(0.0,0.0); 
        (C[8] *> O[2])=(0.0,0.0); 
        (C[8] *> O[3])=(0.0,0.0); 
        (C[8] *> O[4])=(0.0,0.0); 
        (C[8] *> O[5])=(0.0,0.0); 
        (C[8] *> O[6])=(0.0,0.0); 
        (C[8] *> O[7])=(0.0,0.0); 
        (C[8] *> O[8])=(0.0,0.0); 
        (C[8] *> O[9])=(0.0,0.0); 
        (C[8] *> O[10])=(0.0,0.0); 
        (C[8] *> O[11])=(0.0,0.0); 
        (C[8] *> O[12])=(0.0,0.0); 
        (C[8] *> O[13])=(0.0,0.0); 
        (C[8] *> O[14])=(0.0,0.0); 
        (C[8] *> O[15])=(0.0,0.0); 
        (C[8] *> O[16])=(0.0,0.0); 
        (C[8] *> O[17])=(0.0,0.0); 
        (C[8] *> O[18])=(0.0,0.0); 
        (C[8] *> O[19])=(0.0,0.0); 
        (C[8] *> O[20])=(0.0,0.0); 
        (C[8] *> O[21])=(0.0,0.0); 
        (C[8] *> O[22])=(0.0,0.0); 
        (C[8] *> O[23])=(0.0,0.0); 
        (C[8] *> O[24])=(0.0,0.0); 
        (C[8] *> O[25])=(0.0,0.0); 
        (C[8] *> O[26])=(0.0,0.0); 
        (C[8] *> O[27])=(0.0,0.0); 
        (C[8] *> O[28])=(0.0,0.0); 
        (C[8] *> O[29])=(0.0,0.0); 
        (C[8] *> O[30])=(0.0,0.0); 
        (C[8] *> O[31])=(0.0,0.0); 
        (C[9] *> O[0])=(0.0,0.0); 
        (C[9] *> O[1])=(0.0,0.0); 
        (C[9] *> O[2])=(0.0,0.0); 
        (C[9] *> O[3])=(0.0,0.0); 
        (C[9] *> O[4])=(0.0,0.0); 
        (C[9] *> O[5])=(0.0,0.0); 
        (C[9] *> O[6])=(0.0,0.0); 
        (C[9] *> O[7])=(0.0,0.0); 
        (C[9] *> O[8])=(0.0,0.0); 
        (C[9] *> O[9])=(0.0,0.0); 
        (C[9] *> O[10])=(0.0,0.0); 
        (C[9] *> O[11])=(0.0,0.0); 
        (C[9] *> O[12])=(0.0,0.0); 
        (C[9] *> O[13])=(0.0,0.0); 
        (C[9] *> O[14])=(0.0,0.0); 
        (C[9] *> O[15])=(0.0,0.0); 
        (C[9] *> O[16])=(0.0,0.0); 
        (C[9] *> O[17])=(0.0,0.0); 
        (C[9] *> O[18])=(0.0,0.0); 
        (C[9] *> O[19])=(0.0,0.0); 
        (C[9] *> O[20])=(0.0,0.0); 
        (C[9] *> O[21])=(0.0,0.0); 
        (C[9] *> O[22])=(0.0,0.0); 
        (C[9] *> O[23])=(0.0,0.0); 
        (C[9] *> O[24])=(0.0,0.0); 
        (C[9] *> O[25])=(0.0,0.0); 
        (C[9] *> O[26])=(0.0,0.0); 
        (C[9] *> O[27])=(0.0,0.0); 
        (C[9] *> O[28])=(0.0,0.0); 
        (C[9] *> O[29])=(0.0,0.0); 
        (C[9] *> O[30])=(0.0,0.0); 
        (C[9] *> O[31])=(0.0,0.0); 
        (C[10] *> O[0])=(0.0,0.0); 
        (C[10] *> O[1])=(0.0,0.0); 
        (C[10] *> O[2])=(0.0,0.0); 
        (C[10] *> O[3])=(0.0,0.0); 
        (C[10] *> O[4])=(0.0,0.0); 
        (C[10] *> O[5])=(0.0,0.0); 
        (C[10] *> O[6])=(0.0,0.0); 
        (C[10] *> O[7])=(0.0,0.0); 
        (C[10] *> O[8])=(0.0,0.0); 
        (C[10] *> O[9])=(0.0,0.0); 
        (C[10] *> O[10])=(0.0,0.0); 
        (C[10] *> O[11])=(0.0,0.0); 
        (C[10] *> O[12])=(0.0,0.0); 
        (C[10] *> O[13])=(0.0,0.0); 
        (C[10] *> O[14])=(0.0,0.0); 
        (C[10] *> O[15])=(0.0,0.0); 
        (C[10] *> O[16])=(0.0,0.0); 
        (C[10] *> O[17])=(0.0,0.0); 
        (C[10] *> O[18])=(0.0,0.0); 
        (C[10] *> O[19])=(0.0,0.0); 
        (C[10] *> O[20])=(0.0,0.0); 
        (C[10] *> O[21])=(0.0,0.0); 
        (C[10] *> O[22])=(0.0,0.0); 
        (C[10] *> O[23])=(0.0,0.0); 
        (C[10] *> O[24])=(0.0,0.0); 
        (C[10] *> O[25])=(0.0,0.0); 
        (C[10] *> O[26])=(0.0,0.0); 
        (C[10] *> O[27])=(0.0,0.0); 
        (C[10] *> O[28])=(0.0,0.0); 
        (C[10] *> O[29])=(0.0,0.0); 
        (C[10] *> O[30])=(0.0,0.0); 
        (C[10] *> O[31])=(0.0,0.0); 
        (C[11] *> O[0])=(0.0,0.0); 
        (C[11] *> O[1])=(0.0,0.0); 
        (C[11] *> O[2])=(0.0,0.0); 
        (C[11] *> O[3])=(0.0,0.0); 
        (C[11] *> O[4])=(0.0,0.0); 
        (C[11] *> O[5])=(0.0,0.0); 
        (C[11] *> O[6])=(0.0,0.0); 
        (C[11] *> O[7])=(0.0,0.0); 
        (C[11] *> O[8])=(0.0,0.0); 
        (C[11] *> O[9])=(0.0,0.0); 
        (C[11] *> O[10])=(0.0,0.0); 
        (C[11] *> O[11])=(0.0,0.0); 
        (C[11] *> O[12])=(0.0,0.0); 
        (C[11] *> O[13])=(0.0,0.0); 
        (C[11] *> O[14])=(0.0,0.0); 
        (C[11] *> O[15])=(0.0,0.0); 
        (C[11] *> O[16])=(0.0,0.0); 
        (C[11] *> O[17])=(0.0,0.0); 
        (C[11] *> O[18])=(0.0,0.0); 
        (C[11] *> O[19])=(0.0,0.0); 
        (C[11] *> O[20])=(0.0,0.0); 
        (C[11] *> O[21])=(0.0,0.0); 
        (C[11] *> O[22])=(0.0,0.0); 
        (C[11] *> O[23])=(0.0,0.0); 
        (C[11] *> O[24])=(0.0,0.0); 
        (C[11] *> O[25])=(0.0,0.0); 
        (C[11] *> O[26])=(0.0,0.0); 
        (C[11] *> O[27])=(0.0,0.0); 
        (C[11] *> O[28])=(0.0,0.0); 
        (C[11] *> O[29])=(0.0,0.0); 
        (C[11] *> O[30])=(0.0,0.0); 
        (C[11] *> O[31])=(0.0,0.0); 
        (C[12] *> O[0])=(0.0,0.0); 
        (C[12] *> O[1])=(0.0,0.0); 
        (C[12] *> O[2])=(0.0,0.0); 
        (C[12] *> O[3])=(0.0,0.0); 
        (C[12] *> O[4])=(0.0,0.0); 
        (C[12] *> O[5])=(0.0,0.0); 
        (C[12] *> O[6])=(0.0,0.0); 
        (C[12] *> O[7])=(0.0,0.0); 
        (C[12] *> O[8])=(0.0,0.0); 
        (C[12] *> O[9])=(0.0,0.0); 
        (C[12] *> O[10])=(0.0,0.0); 
        (C[12] *> O[11])=(0.0,0.0); 
        (C[12] *> O[12])=(0.0,0.0); 
        (C[12] *> O[13])=(0.0,0.0); 
        (C[12] *> O[14])=(0.0,0.0); 
        (C[12] *> O[15])=(0.0,0.0); 
        (C[12] *> O[16])=(0.0,0.0); 
        (C[12] *> O[17])=(0.0,0.0); 
        (C[12] *> O[18])=(0.0,0.0); 
        (C[12] *> O[19])=(0.0,0.0); 
        (C[12] *> O[20])=(0.0,0.0); 
        (C[12] *> O[21])=(0.0,0.0); 
        (C[12] *> O[22])=(0.0,0.0); 
        (C[12] *> O[23])=(0.0,0.0); 
        (C[12] *> O[24])=(0.0,0.0); 
        (C[12] *> O[25])=(0.0,0.0); 
        (C[12] *> O[26])=(0.0,0.0); 
        (C[12] *> O[27])=(0.0,0.0); 
        (C[12] *> O[28])=(0.0,0.0); 
        (C[12] *> O[29])=(0.0,0.0); 
        (C[12] *> O[30])=(0.0,0.0); 
        (C[12] *> O[31])=(0.0,0.0); 
        (C[13] *> O[0])=(0.0,0.0); 
        (C[13] *> O[1])=(0.0,0.0); 
        (C[13] *> O[2])=(0.0,0.0); 
        (C[13] *> O[3])=(0.0,0.0); 
        (C[13] *> O[4])=(0.0,0.0); 
        (C[13] *> O[5])=(0.0,0.0); 
        (C[13] *> O[6])=(0.0,0.0); 
        (C[13] *> O[7])=(0.0,0.0); 
        (C[13] *> O[8])=(0.0,0.0); 
        (C[13] *> O[9])=(0.0,0.0); 
        (C[13] *> O[10])=(0.0,0.0); 
        (C[13] *> O[11])=(0.0,0.0); 
        (C[13] *> O[12])=(0.0,0.0); 
        (C[13] *> O[13])=(0.0,0.0); 
        (C[13] *> O[14])=(0.0,0.0); 
        (C[13] *> O[15])=(0.0,0.0); 
        (C[13] *> O[16])=(0.0,0.0); 
        (C[13] *> O[17])=(0.0,0.0); 
        (C[13] *> O[18])=(0.0,0.0); 
        (C[13] *> O[19])=(0.0,0.0); 
        (C[13] *> O[20])=(0.0,0.0); 
        (C[13] *> O[21])=(0.0,0.0); 
        (C[13] *> O[22])=(0.0,0.0); 
        (C[13] *> O[23])=(0.0,0.0); 
        (C[13] *> O[24])=(0.0,0.0); 
        (C[13] *> O[25])=(0.0,0.0); 
        (C[13] *> O[26])=(0.0,0.0); 
        (C[13] *> O[27])=(0.0,0.0); 
        (C[13] *> O[28])=(0.0,0.0); 
        (C[13] *> O[29])=(0.0,0.0); 
        (C[13] *> O[30])=(0.0,0.0); 
        (C[13] *> O[31])=(0.0,0.0); 
        (C[14] *> O[0])=(0.0,0.0); 
        (C[14] *> O[1])=(0.0,0.0); 
        (C[14] *> O[2])=(0.0,0.0); 
        (C[14] *> O[3])=(0.0,0.0); 
        (C[14] *> O[4])=(0.0,0.0); 
        (C[14] *> O[5])=(0.0,0.0); 
        (C[14] *> O[6])=(0.0,0.0); 
        (C[14] *> O[7])=(0.0,0.0); 
        (C[14] *> O[8])=(0.0,0.0); 
        (C[14] *> O[9])=(0.0,0.0); 
        (C[14] *> O[10])=(0.0,0.0); 
        (C[14] *> O[11])=(0.0,0.0); 
        (C[14] *> O[12])=(0.0,0.0); 
        (C[14] *> O[13])=(0.0,0.0); 
        (C[14] *> O[14])=(0.0,0.0); 
        (C[14] *> O[15])=(0.0,0.0); 
        (C[14] *> O[16])=(0.0,0.0); 
        (C[14] *> O[17])=(0.0,0.0); 
        (C[14] *> O[18])=(0.0,0.0); 
        (C[14] *> O[19])=(0.0,0.0); 
        (C[14] *> O[20])=(0.0,0.0); 
        (C[14] *> O[21])=(0.0,0.0); 
        (C[14] *> O[22])=(0.0,0.0); 
        (C[14] *> O[23])=(0.0,0.0); 
        (C[14] *> O[24])=(0.0,0.0); 
        (C[14] *> O[25])=(0.0,0.0); 
        (C[14] *> O[26])=(0.0,0.0); 
        (C[14] *> O[27])=(0.0,0.0); 
        (C[14] *> O[28])=(0.0,0.0); 
        (C[14] *> O[29])=(0.0,0.0); 
        (C[14] *> O[30])=(0.0,0.0); 
        (C[14] *> O[31])=(0.0,0.0); 
        (C[15] *> O[0])=(0.0,0.0); 
        (C[15] *> O[1])=(0.0,0.0); 
        (C[15] *> O[2])=(0.0,0.0); 
        (C[15] *> O[3])=(0.0,0.0); 
        (C[15] *> O[4])=(0.0,0.0); 
        (C[15] *> O[5])=(0.0,0.0); 
        (C[15] *> O[6])=(0.0,0.0); 
        (C[15] *> O[7])=(0.0,0.0); 
        (C[15] *> O[8])=(0.0,0.0); 
        (C[15] *> O[9])=(0.0,0.0); 
        (C[15] *> O[10])=(0.0,0.0); 
        (C[15] *> O[11])=(0.0,0.0); 
        (C[15] *> O[12])=(0.0,0.0); 
        (C[15] *> O[13])=(0.0,0.0); 
        (C[15] *> O[14])=(0.0,0.0); 
        (C[15] *> O[15])=(0.0,0.0); 
        (C[15] *> O[16])=(0.0,0.0); 
        (C[15] *> O[17])=(0.0,0.0); 
        (C[15] *> O[18])=(0.0,0.0); 
        (C[15] *> O[19])=(0.0,0.0); 
        (C[15] *> O[20])=(0.0,0.0); 
        (C[15] *> O[21])=(0.0,0.0); 
        (C[15] *> O[22])=(0.0,0.0); 
        (C[15] *> O[23])=(0.0,0.0); 
        (C[15] *> O[24])=(0.0,0.0); 
        (C[15] *> O[25])=(0.0,0.0); 
        (C[15] *> O[26])=(0.0,0.0); 
        (C[15] *> O[27])=(0.0,0.0); 
        (C[15] *> O[28])=(0.0,0.0); 
        (C[15] *> O[29])=(0.0,0.0); 
        (C[15] *> O[30])=(0.0,0.0); 
        (C[15] *> O[31])=(0.0,0.0); 
        (D[0] *> O[0])=(0.0,0.0); 
        (D[0] *> O[1])=(0.0,0.0); 
        (D[0] *> O[2])=(0.0,0.0); 
        (D[0] *> O[3])=(0.0,0.0); 
        (D[0] *> O[4])=(0.0,0.0); 
        (D[0] *> O[5])=(0.0,0.0); 
        (D[0] *> O[6])=(0.0,0.0); 
        (D[0] *> O[7])=(0.0,0.0); 
        (D[0] *> O[8])=(0.0,0.0); 
        (D[0] *> O[9])=(0.0,0.0); 
        (D[0] *> O[10])=(0.0,0.0); 
        (D[0] *> O[11])=(0.0,0.0); 
        (D[0] *> O[12])=(0.0,0.0); 
        (D[0] *> O[13])=(0.0,0.0); 
        (D[0] *> O[14])=(0.0,0.0); 
        (D[0] *> O[15])=(0.0,0.0); 
        (D[0] *> O[16])=(0.0,0.0); 
        (D[0] *> O[17])=(0.0,0.0); 
        (D[0] *> O[18])=(0.0,0.0); 
        (D[0] *> O[19])=(0.0,0.0); 
        (D[0] *> O[20])=(0.0,0.0); 
        (D[0] *> O[21])=(0.0,0.0); 
        (D[0] *> O[22])=(0.0,0.0); 
        (D[0] *> O[23])=(0.0,0.0); 
        (D[0] *> O[24])=(0.0,0.0); 
        (D[0] *> O[25])=(0.0,0.0); 
        (D[0] *> O[26])=(0.0,0.0); 
        (D[0] *> O[27])=(0.0,0.0); 
        (D[0] *> O[28])=(0.0,0.0); 
        (D[0] *> O[29])=(0.0,0.0); 
        (D[0] *> O[30])=(0.0,0.0); 
        (D[0] *> O[31])=(0.0,0.0); 
        (D[1] *> O[0])=(0.0,0.0); 
        (D[1] *> O[1])=(0.0,0.0); 
        (D[1] *> O[2])=(0.0,0.0); 
        (D[1] *> O[3])=(0.0,0.0); 
        (D[1] *> O[4])=(0.0,0.0); 
        (D[1] *> O[5])=(0.0,0.0); 
        (D[1] *> O[6])=(0.0,0.0); 
        (D[1] *> O[7])=(0.0,0.0); 
        (D[1] *> O[8])=(0.0,0.0); 
        (D[1] *> O[9])=(0.0,0.0); 
        (D[1] *> O[10])=(0.0,0.0); 
        (D[1] *> O[11])=(0.0,0.0); 
        (D[1] *> O[12])=(0.0,0.0); 
        (D[1] *> O[13])=(0.0,0.0); 
        (D[1] *> O[14])=(0.0,0.0); 
        (D[1] *> O[15])=(0.0,0.0); 
        (D[1] *> O[16])=(0.0,0.0); 
        (D[1] *> O[17])=(0.0,0.0); 
        (D[1] *> O[18])=(0.0,0.0); 
        (D[1] *> O[19])=(0.0,0.0); 
        (D[1] *> O[20])=(0.0,0.0); 
        (D[1] *> O[21])=(0.0,0.0); 
        (D[1] *> O[22])=(0.0,0.0); 
        (D[1] *> O[23])=(0.0,0.0); 
        (D[1] *> O[24])=(0.0,0.0); 
        (D[1] *> O[25])=(0.0,0.0); 
        (D[1] *> O[26])=(0.0,0.0); 
        (D[1] *> O[27])=(0.0,0.0); 
        (D[1] *> O[28])=(0.0,0.0); 
        (D[1] *> O[29])=(0.0,0.0); 
        (D[1] *> O[30])=(0.0,0.0); 
        (D[1] *> O[31])=(0.0,0.0); 
        (D[2] *> O[0])=(0.0,0.0); 
        (D[2] *> O[1])=(0.0,0.0); 
        (D[2] *> O[2])=(0.0,0.0); 
        (D[2] *> O[3])=(0.0,0.0); 
        (D[2] *> O[4])=(0.0,0.0); 
        (D[2] *> O[5])=(0.0,0.0); 
        (D[2] *> O[6])=(0.0,0.0); 
        (D[2] *> O[7])=(0.0,0.0); 
        (D[2] *> O[8])=(0.0,0.0); 
        (D[2] *> O[9])=(0.0,0.0); 
        (D[2] *> O[10])=(0.0,0.0); 
        (D[2] *> O[11])=(0.0,0.0); 
        (D[2] *> O[12])=(0.0,0.0); 
        (D[2] *> O[13])=(0.0,0.0); 
        (D[2] *> O[14])=(0.0,0.0); 
        (D[2] *> O[15])=(0.0,0.0); 
        (D[2] *> O[16])=(0.0,0.0); 
        (D[2] *> O[17])=(0.0,0.0); 
        (D[2] *> O[18])=(0.0,0.0); 
        (D[2] *> O[19])=(0.0,0.0); 
        (D[2] *> O[20])=(0.0,0.0); 
        (D[2] *> O[21])=(0.0,0.0); 
        (D[2] *> O[22])=(0.0,0.0); 
        (D[2] *> O[23])=(0.0,0.0); 
        (D[2] *> O[24])=(0.0,0.0); 
        (D[2] *> O[25])=(0.0,0.0); 
        (D[2] *> O[26])=(0.0,0.0); 
        (D[2] *> O[27])=(0.0,0.0); 
        (D[2] *> O[28])=(0.0,0.0); 
        (D[2] *> O[29])=(0.0,0.0); 
        (D[2] *> O[30])=(0.0,0.0); 
        (D[2] *> O[31])=(0.0,0.0); 
        (D[3] *> O[0])=(0.0,0.0); 
        (D[3] *> O[1])=(0.0,0.0); 
        (D[3] *> O[2])=(0.0,0.0); 
        (D[3] *> O[3])=(0.0,0.0); 
        (D[3] *> O[4])=(0.0,0.0); 
        (D[3] *> O[5])=(0.0,0.0); 
        (D[3] *> O[6])=(0.0,0.0); 
        (D[3] *> O[7])=(0.0,0.0); 
        (D[3] *> O[8])=(0.0,0.0); 
        (D[3] *> O[9])=(0.0,0.0); 
        (D[3] *> O[10])=(0.0,0.0); 
        (D[3] *> O[11])=(0.0,0.0); 
        (D[3] *> O[12])=(0.0,0.0); 
        (D[3] *> O[13])=(0.0,0.0); 
        (D[3] *> O[14])=(0.0,0.0); 
        (D[3] *> O[15])=(0.0,0.0); 
        (D[3] *> O[16])=(0.0,0.0); 
        (D[3] *> O[17])=(0.0,0.0); 
        (D[3] *> O[18])=(0.0,0.0); 
        (D[3] *> O[19])=(0.0,0.0); 
        (D[3] *> O[20])=(0.0,0.0); 
        (D[3] *> O[21])=(0.0,0.0); 
        (D[3] *> O[22])=(0.0,0.0); 
        (D[3] *> O[23])=(0.0,0.0); 
        (D[3] *> O[24])=(0.0,0.0); 
        (D[3] *> O[25])=(0.0,0.0); 
        (D[3] *> O[26])=(0.0,0.0); 
        (D[3] *> O[27])=(0.0,0.0); 
        (D[3] *> O[28])=(0.0,0.0); 
        (D[3] *> O[29])=(0.0,0.0); 
        (D[3] *> O[30])=(0.0,0.0); 
        (D[3] *> O[31])=(0.0,0.0); 
        (D[4] *> O[0])=(0.0,0.0); 
        (D[4] *> O[1])=(0.0,0.0); 
        (D[4] *> O[2])=(0.0,0.0); 
        (D[4] *> O[3])=(0.0,0.0); 
        (D[4] *> O[4])=(0.0,0.0); 
        (D[4] *> O[5])=(0.0,0.0); 
        (D[4] *> O[6])=(0.0,0.0); 
        (D[4] *> O[7])=(0.0,0.0); 
        (D[4] *> O[8])=(0.0,0.0); 
        (D[4] *> O[9])=(0.0,0.0); 
        (D[4] *> O[10])=(0.0,0.0); 
        (D[4] *> O[11])=(0.0,0.0); 
        (D[4] *> O[12])=(0.0,0.0); 
        (D[4] *> O[13])=(0.0,0.0); 
        (D[4] *> O[14])=(0.0,0.0); 
        (D[4] *> O[15])=(0.0,0.0); 
        (D[4] *> O[16])=(0.0,0.0); 
        (D[4] *> O[17])=(0.0,0.0); 
        (D[4] *> O[18])=(0.0,0.0); 
        (D[4] *> O[19])=(0.0,0.0); 
        (D[4] *> O[20])=(0.0,0.0); 
        (D[4] *> O[21])=(0.0,0.0); 
        (D[4] *> O[22])=(0.0,0.0); 
        (D[4] *> O[23])=(0.0,0.0); 
        (D[4] *> O[24])=(0.0,0.0); 
        (D[4] *> O[25])=(0.0,0.0); 
        (D[4] *> O[26])=(0.0,0.0); 
        (D[4] *> O[27])=(0.0,0.0); 
        (D[4] *> O[28])=(0.0,0.0); 
        (D[4] *> O[29])=(0.0,0.0); 
        (D[4] *> O[30])=(0.0,0.0); 
        (D[4] *> O[31])=(0.0,0.0); 
        (D[5] *> O[0])=(0.0,0.0); 
        (D[5] *> O[1])=(0.0,0.0); 
        (D[5] *> O[2])=(0.0,0.0); 
        (D[5] *> O[3])=(0.0,0.0); 
        (D[5] *> O[4])=(0.0,0.0); 
        (D[5] *> O[5])=(0.0,0.0); 
        (D[5] *> O[6])=(0.0,0.0); 
        (D[5] *> O[7])=(0.0,0.0); 
        (D[5] *> O[8])=(0.0,0.0); 
        (D[5] *> O[9])=(0.0,0.0); 
        (D[5] *> O[10])=(0.0,0.0); 
        (D[5] *> O[11])=(0.0,0.0); 
        (D[5] *> O[12])=(0.0,0.0); 
        (D[5] *> O[13])=(0.0,0.0); 
        (D[5] *> O[14])=(0.0,0.0); 
        (D[5] *> O[15])=(0.0,0.0); 
        (D[5] *> O[16])=(0.0,0.0); 
        (D[5] *> O[17])=(0.0,0.0); 
        (D[5] *> O[18])=(0.0,0.0); 
        (D[5] *> O[19])=(0.0,0.0); 
        (D[5] *> O[20])=(0.0,0.0); 
        (D[5] *> O[21])=(0.0,0.0); 
        (D[5] *> O[22])=(0.0,0.0); 
        (D[5] *> O[23])=(0.0,0.0); 
        (D[5] *> O[24])=(0.0,0.0); 
        (D[5] *> O[25])=(0.0,0.0); 
        (D[5] *> O[26])=(0.0,0.0); 
        (D[5] *> O[27])=(0.0,0.0); 
        (D[5] *> O[28])=(0.0,0.0); 
        (D[5] *> O[29])=(0.0,0.0); 
        (D[5] *> O[30])=(0.0,0.0); 
        (D[5] *> O[31])=(0.0,0.0); 
        (D[6] *> O[0])=(0.0,0.0); 
        (D[6] *> O[1])=(0.0,0.0); 
        (D[6] *> O[2])=(0.0,0.0); 
        (D[6] *> O[3])=(0.0,0.0); 
        (D[6] *> O[4])=(0.0,0.0); 
        (D[6] *> O[5])=(0.0,0.0); 
        (D[6] *> O[6])=(0.0,0.0); 
        (D[6] *> O[7])=(0.0,0.0); 
        (D[6] *> O[8])=(0.0,0.0); 
        (D[6] *> O[9])=(0.0,0.0); 
        (D[6] *> O[10])=(0.0,0.0); 
        (D[6] *> O[11])=(0.0,0.0); 
        (D[6] *> O[12])=(0.0,0.0); 
        (D[6] *> O[13])=(0.0,0.0); 
        (D[6] *> O[14])=(0.0,0.0); 
        (D[6] *> O[15])=(0.0,0.0); 
        (D[6] *> O[16])=(0.0,0.0); 
        (D[6] *> O[17])=(0.0,0.0); 
        (D[6] *> O[18])=(0.0,0.0); 
        (D[6] *> O[19])=(0.0,0.0); 
        (D[6] *> O[20])=(0.0,0.0); 
        (D[6] *> O[21])=(0.0,0.0); 
        (D[6] *> O[22])=(0.0,0.0); 
        (D[6] *> O[23])=(0.0,0.0); 
        (D[6] *> O[24])=(0.0,0.0); 
        (D[6] *> O[25])=(0.0,0.0); 
        (D[6] *> O[26])=(0.0,0.0); 
        (D[6] *> O[27])=(0.0,0.0); 
        (D[6] *> O[28])=(0.0,0.0); 
        (D[6] *> O[29])=(0.0,0.0); 
        (D[6] *> O[30])=(0.0,0.0); 
        (D[6] *> O[31])=(0.0,0.0); 
        (D[7] *> O[0])=(0.0,0.0); 
        (D[7] *> O[1])=(0.0,0.0); 
        (D[7] *> O[2])=(0.0,0.0); 
        (D[7] *> O[3])=(0.0,0.0); 
        (D[7] *> O[4])=(0.0,0.0); 
        (D[7] *> O[5])=(0.0,0.0); 
        (D[7] *> O[6])=(0.0,0.0); 
        (D[7] *> O[7])=(0.0,0.0); 
        (D[7] *> O[8])=(0.0,0.0); 
        (D[7] *> O[9])=(0.0,0.0); 
        (D[7] *> O[10])=(0.0,0.0); 
        (D[7] *> O[11])=(0.0,0.0); 
        (D[7] *> O[12])=(0.0,0.0); 
        (D[7] *> O[13])=(0.0,0.0); 
        (D[7] *> O[14])=(0.0,0.0); 
        (D[7] *> O[15])=(0.0,0.0); 
        (D[7] *> O[16])=(0.0,0.0); 
        (D[7] *> O[17])=(0.0,0.0); 
        (D[7] *> O[18])=(0.0,0.0); 
        (D[7] *> O[19])=(0.0,0.0); 
        (D[7] *> O[20])=(0.0,0.0); 
        (D[7] *> O[21])=(0.0,0.0); 
        (D[7] *> O[22])=(0.0,0.0); 
        (D[7] *> O[23])=(0.0,0.0); 
        (D[7] *> O[24])=(0.0,0.0); 
        (D[7] *> O[25])=(0.0,0.0); 
        (D[7] *> O[26])=(0.0,0.0); 
        (D[7] *> O[27])=(0.0,0.0); 
        (D[7] *> O[28])=(0.0,0.0); 
        (D[7] *> O[29])=(0.0,0.0); 
        (D[7] *> O[30])=(0.0,0.0); 
        (D[7] *> O[31])=(0.0,0.0); 
        (D[8] *> O[0])=(0.0,0.0); 
        (D[8] *> O[1])=(0.0,0.0); 
        (D[8] *> O[2])=(0.0,0.0); 
        (D[8] *> O[3])=(0.0,0.0); 
        (D[8] *> O[4])=(0.0,0.0); 
        (D[8] *> O[5])=(0.0,0.0); 
        (D[8] *> O[6])=(0.0,0.0); 
        (D[8] *> O[7])=(0.0,0.0); 
        (D[8] *> O[8])=(0.0,0.0); 
        (D[8] *> O[9])=(0.0,0.0); 
        (D[8] *> O[10])=(0.0,0.0); 
        (D[8] *> O[11])=(0.0,0.0); 
        (D[8] *> O[12])=(0.0,0.0); 
        (D[8] *> O[13])=(0.0,0.0); 
        (D[8] *> O[14])=(0.0,0.0); 
        (D[8] *> O[15])=(0.0,0.0); 
        (D[8] *> O[16])=(0.0,0.0); 
        (D[8] *> O[17])=(0.0,0.0); 
        (D[8] *> O[18])=(0.0,0.0); 
        (D[8] *> O[19])=(0.0,0.0); 
        (D[8] *> O[20])=(0.0,0.0); 
        (D[8] *> O[21])=(0.0,0.0); 
        (D[8] *> O[22])=(0.0,0.0); 
        (D[8] *> O[23])=(0.0,0.0); 
        (D[8] *> O[24])=(0.0,0.0); 
        (D[8] *> O[25])=(0.0,0.0); 
        (D[8] *> O[26])=(0.0,0.0); 
        (D[8] *> O[27])=(0.0,0.0); 
        (D[8] *> O[28])=(0.0,0.0); 
        (D[8] *> O[29])=(0.0,0.0); 
        (D[8] *> O[30])=(0.0,0.0); 
        (D[8] *> O[31])=(0.0,0.0); 
        (D[9] *> O[0])=(0.0,0.0); 
        (D[9] *> O[1])=(0.0,0.0); 
        (D[9] *> O[2])=(0.0,0.0); 
        (D[9] *> O[3])=(0.0,0.0); 
        (D[9] *> O[4])=(0.0,0.0); 
        (D[9] *> O[5])=(0.0,0.0); 
        (D[9] *> O[6])=(0.0,0.0); 
        (D[9] *> O[7])=(0.0,0.0); 
        (D[9] *> O[8])=(0.0,0.0); 
        (D[9] *> O[9])=(0.0,0.0); 
        (D[9] *> O[10])=(0.0,0.0); 
        (D[9] *> O[11])=(0.0,0.0); 
        (D[9] *> O[12])=(0.0,0.0); 
        (D[9] *> O[13])=(0.0,0.0); 
        (D[9] *> O[14])=(0.0,0.0); 
        (D[9] *> O[15])=(0.0,0.0); 
        (D[9] *> O[16])=(0.0,0.0); 
        (D[9] *> O[17])=(0.0,0.0); 
        (D[9] *> O[18])=(0.0,0.0); 
        (D[9] *> O[19])=(0.0,0.0); 
        (D[9] *> O[20])=(0.0,0.0); 
        (D[9] *> O[21])=(0.0,0.0); 
        (D[9] *> O[22])=(0.0,0.0); 
        (D[9] *> O[23])=(0.0,0.0); 
        (D[9] *> O[24])=(0.0,0.0); 
        (D[9] *> O[25])=(0.0,0.0); 
        (D[9] *> O[26])=(0.0,0.0); 
        (D[9] *> O[27])=(0.0,0.0); 
        (D[9] *> O[28])=(0.0,0.0); 
        (D[9] *> O[29])=(0.0,0.0); 
        (D[9] *> O[30])=(0.0,0.0); 
        (D[9] *> O[31])=(0.0,0.0); 
        (D[10] *> O[0])=(0.0,0.0); 
        (D[10] *> O[1])=(0.0,0.0); 
        (D[10] *> O[2])=(0.0,0.0); 
        (D[10] *> O[3])=(0.0,0.0); 
        (D[10] *> O[4])=(0.0,0.0); 
        (D[10] *> O[5])=(0.0,0.0); 
        (D[10] *> O[6])=(0.0,0.0); 
        (D[10] *> O[7])=(0.0,0.0); 
        (D[10] *> O[8])=(0.0,0.0); 
        (D[10] *> O[9])=(0.0,0.0); 
        (D[10] *> O[10])=(0.0,0.0); 
        (D[10] *> O[11])=(0.0,0.0); 
        (D[10] *> O[12])=(0.0,0.0); 
        (D[10] *> O[13])=(0.0,0.0); 
        (D[10] *> O[14])=(0.0,0.0); 
        (D[10] *> O[15])=(0.0,0.0); 
        (D[10] *> O[16])=(0.0,0.0); 
        (D[10] *> O[17])=(0.0,0.0); 
        (D[10] *> O[18])=(0.0,0.0); 
        (D[10] *> O[19])=(0.0,0.0); 
        (D[10] *> O[20])=(0.0,0.0); 
        (D[10] *> O[21])=(0.0,0.0); 
        (D[10] *> O[22])=(0.0,0.0); 
        (D[10] *> O[23])=(0.0,0.0); 
        (D[10] *> O[24])=(0.0,0.0); 
        (D[10] *> O[25])=(0.0,0.0); 
        (D[10] *> O[26])=(0.0,0.0); 
        (D[10] *> O[27])=(0.0,0.0); 
        (D[10] *> O[28])=(0.0,0.0); 
        (D[10] *> O[29])=(0.0,0.0); 
        (D[10] *> O[30])=(0.0,0.0); 
        (D[10] *> O[31])=(0.0,0.0); 
        (D[11] *> O[0])=(0.0,0.0); 
        (D[11] *> O[1])=(0.0,0.0); 
        (D[11] *> O[2])=(0.0,0.0); 
        (D[11] *> O[3])=(0.0,0.0); 
        (D[11] *> O[4])=(0.0,0.0); 
        (D[11] *> O[5])=(0.0,0.0); 
        (D[11] *> O[6])=(0.0,0.0); 
        (D[11] *> O[7])=(0.0,0.0); 
        (D[11] *> O[8])=(0.0,0.0); 
        (D[11] *> O[9])=(0.0,0.0); 
        (D[11] *> O[10])=(0.0,0.0); 
        (D[11] *> O[11])=(0.0,0.0); 
        (D[11] *> O[12])=(0.0,0.0); 
        (D[11] *> O[13])=(0.0,0.0); 
        (D[11] *> O[14])=(0.0,0.0); 
        (D[11] *> O[15])=(0.0,0.0); 
        (D[11] *> O[16])=(0.0,0.0); 
        (D[11] *> O[17])=(0.0,0.0); 
        (D[11] *> O[18])=(0.0,0.0); 
        (D[11] *> O[19])=(0.0,0.0); 
        (D[11] *> O[20])=(0.0,0.0); 
        (D[11] *> O[21])=(0.0,0.0); 
        (D[11] *> O[22])=(0.0,0.0); 
        (D[11] *> O[23])=(0.0,0.0); 
        (D[11] *> O[24])=(0.0,0.0); 
        (D[11] *> O[25])=(0.0,0.0); 
        (D[11] *> O[26])=(0.0,0.0); 
        (D[11] *> O[27])=(0.0,0.0); 
        (D[11] *> O[28])=(0.0,0.0); 
        (D[11] *> O[29])=(0.0,0.0); 
        (D[11] *> O[30])=(0.0,0.0); 
        (D[11] *> O[31])=(0.0,0.0); 
        (D[12] *> O[0])=(0.0,0.0); 
        (D[12] *> O[1])=(0.0,0.0); 
        (D[12] *> O[2])=(0.0,0.0); 
        (D[12] *> O[3])=(0.0,0.0); 
        (D[12] *> O[4])=(0.0,0.0); 
        (D[12] *> O[5])=(0.0,0.0); 
        (D[12] *> O[6])=(0.0,0.0); 
        (D[12] *> O[7])=(0.0,0.0); 
        (D[12] *> O[8])=(0.0,0.0); 
        (D[12] *> O[9])=(0.0,0.0); 
        (D[12] *> O[10])=(0.0,0.0); 
        (D[12] *> O[11])=(0.0,0.0); 
        (D[12] *> O[12])=(0.0,0.0); 
        (D[12] *> O[13])=(0.0,0.0); 
        (D[12] *> O[14])=(0.0,0.0); 
        (D[12] *> O[15])=(0.0,0.0); 
        (D[12] *> O[16])=(0.0,0.0); 
        (D[12] *> O[17])=(0.0,0.0); 
        (D[12] *> O[18])=(0.0,0.0); 
        (D[12] *> O[19])=(0.0,0.0); 
        (D[12] *> O[20])=(0.0,0.0); 
        (D[12] *> O[21])=(0.0,0.0); 
        (D[12] *> O[22])=(0.0,0.0); 
        (D[12] *> O[23])=(0.0,0.0); 
        (D[12] *> O[24])=(0.0,0.0); 
        (D[12] *> O[25])=(0.0,0.0); 
        (D[12] *> O[26])=(0.0,0.0); 
        (D[12] *> O[27])=(0.0,0.0); 
        (D[12] *> O[28])=(0.0,0.0); 
        (D[12] *> O[29])=(0.0,0.0); 
        (D[12] *> O[30])=(0.0,0.0); 
        (D[12] *> O[31])=(0.0,0.0); 
        (D[13] *> O[0])=(0.0,0.0); 
        (D[13] *> O[1])=(0.0,0.0); 
        (D[13] *> O[2])=(0.0,0.0); 
        (D[13] *> O[3])=(0.0,0.0); 
        (D[13] *> O[4])=(0.0,0.0); 
        (D[13] *> O[5])=(0.0,0.0); 
        (D[13] *> O[6])=(0.0,0.0); 
        (D[13] *> O[7])=(0.0,0.0); 
        (D[13] *> O[8])=(0.0,0.0); 
        (D[13] *> O[9])=(0.0,0.0); 
        (D[13] *> O[10])=(0.0,0.0); 
        (D[13] *> O[11])=(0.0,0.0); 
        (D[13] *> O[12])=(0.0,0.0); 
        (D[13] *> O[13])=(0.0,0.0); 
        (D[13] *> O[14])=(0.0,0.0); 
        (D[13] *> O[15])=(0.0,0.0); 
        (D[13] *> O[16])=(0.0,0.0); 
        (D[13] *> O[17])=(0.0,0.0); 
        (D[13] *> O[18])=(0.0,0.0); 
        (D[13] *> O[19])=(0.0,0.0); 
        (D[13] *> O[20])=(0.0,0.0); 
        (D[13] *> O[21])=(0.0,0.0); 
        (D[13] *> O[22])=(0.0,0.0); 
        (D[13] *> O[23])=(0.0,0.0); 
        (D[13] *> O[24])=(0.0,0.0); 
        (D[13] *> O[25])=(0.0,0.0); 
        (D[13] *> O[26])=(0.0,0.0); 
        (D[13] *> O[27])=(0.0,0.0); 
        (D[13] *> O[28])=(0.0,0.0); 
        (D[13] *> O[29])=(0.0,0.0); 
        (D[13] *> O[30])=(0.0,0.0); 
        (D[13] *> O[31])=(0.0,0.0); 
        (D[14] *> O[0])=(0.0,0.0); 
        (D[14] *> O[1])=(0.0,0.0); 
        (D[14] *> O[2])=(0.0,0.0); 
        (D[14] *> O[3])=(0.0,0.0); 
        (D[14] *> O[4])=(0.0,0.0); 
        (D[14] *> O[5])=(0.0,0.0); 
        (D[14] *> O[6])=(0.0,0.0); 
        (D[14] *> O[7])=(0.0,0.0); 
        (D[14] *> O[8])=(0.0,0.0); 
        (D[14] *> O[9])=(0.0,0.0); 
        (D[14] *> O[10])=(0.0,0.0); 
        (D[14] *> O[11])=(0.0,0.0); 
        (D[14] *> O[12])=(0.0,0.0); 
        (D[14] *> O[13])=(0.0,0.0); 
        (D[14] *> O[14])=(0.0,0.0); 
        (D[14] *> O[15])=(0.0,0.0); 
        (D[14] *> O[16])=(0.0,0.0); 
        (D[14] *> O[17])=(0.0,0.0); 
        (D[14] *> O[18])=(0.0,0.0); 
        (D[14] *> O[19])=(0.0,0.0); 
        (D[14] *> O[20])=(0.0,0.0); 
        (D[14] *> O[21])=(0.0,0.0); 
        (D[14] *> O[22])=(0.0,0.0); 
        (D[14] *> O[23])=(0.0,0.0); 
        (D[14] *> O[24])=(0.0,0.0); 
        (D[14] *> O[25])=(0.0,0.0); 
        (D[14] *> O[26])=(0.0,0.0); 
        (D[14] *> O[27])=(0.0,0.0); 
        (D[14] *> O[28])=(0.0,0.0); 
        (D[14] *> O[29])=(0.0,0.0); 
        (D[14] *> O[30])=(0.0,0.0); 
        (D[14] *> O[31])=(0.0,0.0); 
        (D[15] *> O[0])=(0.0,0.0); 
        (D[15] *> O[1])=(0.0,0.0); 
        (D[15] *> O[2])=(0.0,0.0); 
        (D[15] *> O[3])=(0.0,0.0); 
        (D[15] *> O[4])=(0.0,0.0); 
        (D[15] *> O[5])=(0.0,0.0); 
        (D[15] *> O[6])=(0.0,0.0); 
        (D[15] *> O[7])=(0.0,0.0); 
        (D[15] *> O[8])=(0.0,0.0); 
        (D[15] *> O[9])=(0.0,0.0); 
        (D[15] *> O[10])=(0.0,0.0); 
        (D[15] *> O[11])=(0.0,0.0); 
        (D[15] *> O[12])=(0.0,0.0); 
        (D[15] *> O[13])=(0.0,0.0); 
        (D[15] *> O[14])=(0.0,0.0); 
        (D[15] *> O[15])=(0.0,0.0); 
        (D[15] *> O[16])=(0.0,0.0); 
        (D[15] *> O[17])=(0.0,0.0); 
        (D[15] *> O[18])=(0.0,0.0); 
        (D[15] *> O[19])=(0.0,0.0); 
        (D[15] *> O[20])=(0.0,0.0); 
        (D[15] *> O[21])=(0.0,0.0); 
        (D[15] *> O[22])=(0.0,0.0); 
        (D[15] *> O[23])=(0.0,0.0); 
        (D[15] *> O[24])=(0.0,0.0); 
        (D[15] *> O[25])=(0.0,0.0); 
        (D[15] *> O[26])=(0.0,0.0); 
        (D[15] *> O[27])=(0.0,0.0); 
        (D[15] *> O[28])=(0.0,0.0); 
        (D[15] *> O[29])=(0.0,0.0); 
        (D[15] *> O[30])=(0.0,0.0); 
        (D[15] *> O[31])=(0.0,0.0); 
        (IRSTBOT *> O[0])=(0.0,0.0); 
        (IRSTBOT *> O[1])=(0.0,0.0); 
        (IRSTBOT *> O[2])=(0.0,0.0); 
        (IRSTBOT *> O[3])=(0.0,0.0); 
        (IRSTBOT *> O[4])=(0.0,0.0); 
        (IRSTBOT *> O[5])=(0.0,0.0); 
        (IRSTBOT *> O[6])=(0.0,0.0); 
        (IRSTBOT *> O[7])=(0.0,0.0); 
        (IRSTBOT *> O[8])=(0.0,0.0); 
        (IRSTBOT *> O[9])=(0.0,0.0); 
        (IRSTBOT *> O[10])=(0.0,0.0); 
        (IRSTBOT *> O[11])=(0.0,0.0); 
        (IRSTBOT *> O[12])=(0.0,0.0); 
        (IRSTBOT *> O[13])=(0.0,0.0); 
        (IRSTBOT *> O[14])=(0.0,0.0); 
        (IRSTBOT *> O[15])=(0.0,0.0); 
        (IRSTBOT *> O[16])=(0.0,0.0); 
        (IRSTBOT *> O[17])=(0.0,0.0); 
        (IRSTBOT *> O[18])=(0.0,0.0); 
        (IRSTBOT *> O[19])=(0.0,0.0); 
        (IRSTBOT *> O[20])=(0.0,0.0); 
        (IRSTBOT *> O[21])=(0.0,0.0); 
        (IRSTBOT *> O[22])=(0.0,0.0); 
        (IRSTBOT *> O[23])=(0.0,0.0); 
        (IRSTBOT *> O[24])=(0.0,0.0); 
        (IRSTBOT *> O[25])=(0.0,0.0); 
        (IRSTBOT *> O[26])=(0.0,0.0); 
        (IRSTBOT *> O[27])=(0.0,0.0); 
        (IRSTBOT *> O[28])=(0.0,0.0); 
        (IRSTBOT *> O[29])=(0.0,0.0); 
        (IRSTBOT *> O[30])=(0.0,0.0); 
        (IRSTBOT *> O[31])=(0.0,0.0); 
        (ORSTBOT *> O[0])=(0.0,0.0); 
        (ORSTBOT *> O[1])=(0.0,0.0); 
        (ORSTBOT *> O[2])=(0.0,0.0); 
        (ORSTBOT *> O[3])=(0.0,0.0); 
        (ORSTBOT *> O[4])=(0.0,0.0); 
        (ORSTBOT *> O[5])=(0.0,0.0); 
        (ORSTBOT *> O[6])=(0.0,0.0); 
        (ORSTBOT *> O[7])=(0.0,0.0); 
        (ORSTBOT *> O[8])=(0.0,0.0); 
        (ORSTBOT *> O[9])=(0.0,0.0); 
        (ORSTBOT *> O[10])=(0.0,0.0); 
        (ORSTBOT *> O[11])=(0.0,0.0); 
        (ORSTBOT *> O[12])=(0.0,0.0); 
        (ORSTBOT *> O[13])=(0.0,0.0); 
        (ORSTBOT *> O[14])=(0.0,0.0); 
        (ORSTBOT *> O[15])=(0.0,0.0); 
        (ORSTBOT *> O[16])=(0.0,0.0); 
        (ORSTBOT *> O[17])=(0.0,0.0); 
        (ORSTBOT *> O[18])=(0.0,0.0); 
        (ORSTBOT *> O[19])=(0.0,0.0); 
        (ORSTBOT *> O[20])=(0.0,0.0); 
        (ORSTBOT *> O[21])=(0.0,0.0); 
        (ORSTBOT *> O[22])=(0.0,0.0); 
        (ORSTBOT *> O[23])=(0.0,0.0); 
        (ORSTBOT *> O[24])=(0.0,0.0); 
        (ORSTBOT *> O[25])=(0.0,0.0); 
        (ORSTBOT *> O[26])=(0.0,0.0); 
        (ORSTBOT *> O[27])=(0.0,0.0); 
        (ORSTBOT *> O[28])=(0.0,0.0); 
        (ORSTBOT *> O[29])=(0.0,0.0); 
        (ORSTBOT *> O[30])=(0.0,0.0); 
        (ORSTBOT *> O[31])=(0.0,0.0); 
        (ORSTTOP *> O[0])=(0.0,0.0); 
        (ORSTTOP *> O[1])=(0.0,0.0); 
        (ORSTTOP *> O[2])=(0.0,0.0); 
        (ORSTTOP *> O[3])=(0.0,0.0); 
        (ORSTTOP *> O[4])=(0.0,0.0); 
        (ORSTTOP *> O[5])=(0.0,0.0); 
        (ORSTTOP *> O[6])=(0.0,0.0); 
        (ORSTTOP *> O[7])=(0.0,0.0); 
        (ORSTTOP *> O[8])=(0.0,0.0); 
        (ORSTTOP *> O[9])=(0.0,0.0); 
        (ORSTTOP *> O[10])=(0.0,0.0); 
        (ORSTTOP *> O[11])=(0.0,0.0); 
        (ORSTTOP *> O[12])=(0.0,0.0); 
        (ORSTTOP *> O[13])=(0.0,0.0); 
        (ORSTTOP *> O[14])=(0.0,0.0); 
        (ORSTTOP *> O[15])=(0.0,0.0); 
        (ORSTTOP *> O[16])=(0.0,0.0); 
        (ORSTTOP *> O[17])=(0.0,0.0); 
        (ORSTTOP *> O[18])=(0.0,0.0); 
        (ORSTTOP *> O[19])=(0.0,0.0); 
        (ORSTTOP *> O[20])=(0.0,0.0); 
        (ORSTTOP *> O[21])=(0.0,0.0); 
        (ORSTTOP *> O[22])=(0.0,0.0); 
        (ORSTTOP *> O[23])=(0.0,0.0); 
        (ORSTTOP *> O[24])=(0.0,0.0); 
        (ORSTTOP *> O[25])=(0.0,0.0); 
        (ORSTTOP *> O[26])=(0.0,0.0); 
        (ORSTTOP *> O[27])=(0.0,0.0); 
        (ORSTTOP *> O[28])=(0.0,0.0); 
        (ORSTTOP *> O[29])=(0.0,0.0); 
        (ORSTTOP *> O[30])=(0.0,0.0); 
        (ORSTTOP *> O[31])=(0.0,0.0); 
        (OLOADTOP *> O[0])=(0.0,0.0); 
        (OLOADTOP *> O[1])=(0.0,0.0); 
        (OLOADTOP *> O[2])=(0.0,0.0); 
        (OLOADTOP *> O[3])=(0.0,0.0); 
        (OLOADTOP *> O[4])=(0.0,0.0); 
        (OLOADTOP *> O[5])=(0.0,0.0); 
        (OLOADTOP *> O[6])=(0.0,0.0); 
        (OLOADTOP *> O[7])=(0.0,0.0); 
        (OLOADTOP *> O[8])=(0.0,0.0); 
        (OLOADTOP *> O[9])=(0.0,0.0); 
        (OLOADTOP *> O[10])=(0.0,0.0); 
        (OLOADTOP *> O[11])=(0.0,0.0); 
        (OLOADTOP *> O[12])=(0.0,0.0); 
        (OLOADTOP *> O[13])=(0.0,0.0); 
        (OLOADTOP *> O[14])=(0.0,0.0); 
        (OLOADTOP *> O[15])=(0.0,0.0); 
        (OLOADTOP *> O[16])=(0.0,0.0); 
        (OLOADTOP *> O[17])=(0.0,0.0); 
        (OLOADTOP *> O[18])=(0.0,0.0); 
        (OLOADTOP *> O[19])=(0.0,0.0); 
        (OLOADTOP *> O[20])=(0.0,0.0); 
        (OLOADTOP *> O[21])=(0.0,0.0); 
        (OLOADTOP *> O[22])=(0.0,0.0); 
        (OLOADTOP *> O[23])=(0.0,0.0); 
        (OLOADTOP *> O[24])=(0.0,0.0); 
        (OLOADTOP *> O[25])=(0.0,0.0); 
        (OLOADTOP *> O[26])=(0.0,0.0); 
        (OLOADTOP *> O[27])=(0.0,0.0); 
        (OLOADTOP *> O[28])=(0.0,0.0); 
        (OLOADTOP *> O[29])=(0.0,0.0); 
        (OLOADTOP *> O[30])=(0.0,0.0); 
        (OLOADTOP *> O[31])=(0.0,0.0); 
        (OLOADBOT *> O[0])=(0.0,0.0); 
        (OLOADBOT *> O[1])=(0.0,0.0); 
        (OLOADBOT *> O[2])=(0.0,0.0); 
        (OLOADBOT *> O[3])=(0.0,0.0); 
        (OLOADBOT *> O[4])=(0.0,0.0); 
        (OLOADBOT *> O[5])=(0.0,0.0); 
        (OLOADBOT *> O[6])=(0.0,0.0); 
        (OLOADBOT *> O[7])=(0.0,0.0); 
        (OLOADBOT *> O[8])=(0.0,0.0); 
        (OLOADBOT *> O[9])=(0.0,0.0); 
        (OLOADBOT *> O[10])=(0.0,0.0); 
        (OLOADBOT *> O[11])=(0.0,0.0); 
        (OLOADBOT *> O[12])=(0.0,0.0); 
        (OLOADBOT *> O[13])=(0.0,0.0); 
        (OLOADBOT *> O[14])=(0.0,0.0); 
        (OLOADBOT *> O[15])=(0.0,0.0); 
        (OLOADBOT *> O[16])=(0.0,0.0); 
        (OLOADBOT *> O[17])=(0.0,0.0); 
        (OLOADBOT *> O[18])=(0.0,0.0); 
        (OLOADBOT *> O[19])=(0.0,0.0); 
        (OLOADBOT *> O[20])=(0.0,0.0); 
        (OLOADBOT *> O[21])=(0.0,0.0); 
        (OLOADBOT *> O[22])=(0.0,0.0); 
        (OLOADBOT *> O[23])=(0.0,0.0); 
        (OLOADBOT *> O[24])=(0.0,0.0); 
        (OLOADBOT *> O[25])=(0.0,0.0); 
        (OLOADBOT *> O[26])=(0.0,0.0); 
        (OLOADBOT *> O[27])=(0.0,0.0); 
        (OLOADBOT *> O[28])=(0.0,0.0); 
        (OLOADBOT *> O[29])=(0.0,0.0); 
        (OLOADBOT *> O[30])=(0.0,0.0); 
        (OLOADBOT *> O[31])=(0.0,0.0); 
      (OLOADTOP *> CO)=(0.0,0.0);
      (OLOADBOT *> CO)=(0.0,0.0);
      (OLOADTOP *> ACCUMCO)=(0.0,0.0);
      (OLOADBOT *> ACCUMCO)=(0.0,0.0);
        (ADDSUBTOP *> O[0])=(0.0,0.0); 
        (ADDSUBTOP *> O[1])=(0.0,0.0); 
        (ADDSUBTOP *> O[2])=(0.0,0.0); 
        (ADDSUBTOP *> O[3])=(0.0,0.0); 
        (ADDSUBTOP *> O[4])=(0.0,0.0); 
        (ADDSUBTOP *> O[5])=(0.0,0.0); 
        (ADDSUBTOP *> O[6])=(0.0,0.0); 
        (ADDSUBTOP *> O[7])=(0.0,0.0); 
        (ADDSUBTOP *> O[8])=(0.0,0.0); 
        (ADDSUBTOP *> O[9])=(0.0,0.0); 
        (ADDSUBTOP *> O[10])=(0.0,0.0); 
        (ADDSUBTOP *> O[11])=(0.0,0.0); 
        (ADDSUBTOP *> O[12])=(0.0,0.0); 
        (ADDSUBTOP *> O[13])=(0.0,0.0); 
        (ADDSUBTOP *> O[14])=(0.0,0.0); 
        (ADDSUBTOP *> O[15])=(0.0,0.0); 
        (ADDSUBTOP *> O[16])=(0.0,0.0); 
        (ADDSUBTOP *> O[17])=(0.0,0.0); 
        (ADDSUBTOP *> O[18])=(0.0,0.0); 
        (ADDSUBTOP *> O[19])=(0.0,0.0); 
        (ADDSUBTOP *> O[20])=(0.0,0.0); 
        (ADDSUBTOP *> O[21])=(0.0,0.0); 
        (ADDSUBTOP *> O[22])=(0.0,0.0); 
        (ADDSUBTOP *> O[23])=(0.0,0.0); 
        (ADDSUBTOP *> O[24])=(0.0,0.0); 
        (ADDSUBTOP *> O[25])=(0.0,0.0); 
        (ADDSUBTOP *> O[26])=(0.0,0.0); 
        (ADDSUBTOP *> O[27])=(0.0,0.0); 
        (ADDSUBTOP *> O[28])=(0.0,0.0); 
        (ADDSUBTOP *> O[29])=(0.0,0.0); 
        (ADDSUBTOP *> O[30])=(0.0,0.0); 
        (ADDSUBTOP *> O[31])=(0.0,0.0); 
        (ADDSUBBOT *> O[0])=(0.0,0.0); 
        (ADDSUBBOT *> O[1])=(0.0,0.0); 
        (ADDSUBBOT *> O[2])=(0.0,0.0); 
        (ADDSUBBOT *> O[3])=(0.0,0.0); 
        (ADDSUBBOT *> O[4])=(0.0,0.0); 
        (ADDSUBBOT *> O[5])=(0.0,0.0); 
        (ADDSUBBOT *> O[6])=(0.0,0.0); 
        (ADDSUBBOT *> O[7])=(0.0,0.0); 
        (ADDSUBBOT *> O[8])=(0.0,0.0); 
        (ADDSUBBOT *> O[9])=(0.0,0.0); 
        (ADDSUBBOT *> O[10])=(0.0,0.0); 
        (ADDSUBBOT *> O[11])=(0.0,0.0); 
        (ADDSUBBOT *> O[12])=(0.0,0.0); 
        (ADDSUBBOT *> O[13])=(0.0,0.0); 
        (ADDSUBBOT *> O[14])=(0.0,0.0); 
        (ADDSUBBOT *> O[15])=(0.0,0.0); 
        (ADDSUBBOT *> O[16])=(0.0,0.0); 
        (ADDSUBBOT *> O[17])=(0.0,0.0); 
        (ADDSUBBOT *> O[18])=(0.0,0.0); 
        (ADDSUBBOT *> O[19])=(0.0,0.0); 
        (ADDSUBBOT *> O[20])=(0.0,0.0); 
        (ADDSUBBOT *> O[21])=(0.0,0.0); 
        (ADDSUBBOT *> O[22])=(0.0,0.0); 
        (ADDSUBBOT *> O[23])=(0.0,0.0); 
        (ADDSUBBOT *> O[24])=(0.0,0.0); 
        (ADDSUBBOT *> O[25])=(0.0,0.0); 
        (ADDSUBBOT *> O[26])=(0.0,0.0); 
        (ADDSUBBOT *> O[27])=(0.0,0.0); 
        (ADDSUBBOT *> O[28])=(0.0,0.0); 
        (ADDSUBBOT *> O[29])=(0.0,0.0); 
        (ADDSUBBOT *> O[30])=(0.0,0.0); 
        (ADDSUBBOT *> O[31])=(0.0,0.0); 
      (ADDSUBTOP *> CO)=(0.0,0.0);
      (ADDSUBBOT *> CO)=(0.0,0.0);
      (ADDSUBTOP *> ACCUMCO)=(0.0,0.0);
      (ADDSUBBOT *> ACCUMCO)=(0.0,0.0);
        (CLK *> O[0])=(0.0,0.0); 
        (CLK *> O[1])=(0.0,0.0); 
        (CLK *> O[2])=(0.0,0.0); 
        (CLK *> O[3])=(0.0,0.0); 
        (CLK *> O[4])=(0.0,0.0); 
        (CLK *> O[5])=(0.0,0.0); 
        (CLK *> O[6])=(0.0,0.0); 
        (CLK *> O[7])=(0.0,0.0); 
        (CLK *> O[8])=(0.0,0.0); 
        (CLK *> O[9])=(0.0,0.0); 
        (CLK *> O[10])=(0.0,0.0); 
        (CLK *> O[11])=(0.0,0.0); 
        (CLK *> O[12])=(0.0,0.0); 
        (CLK *> O[13])=(0.0,0.0); 
        (CLK *> O[14])=(0.0,0.0); 
        (CLK *> O[15])=(0.0,0.0); 
        (CLK *> O[16])=(0.0,0.0); 
        (CLK *> O[17])=(0.0,0.0); 
        (CLK *> O[18])=(0.0,0.0); 
        (CLK *> O[19])=(0.0,0.0); 
        (CLK *> O[20])=(0.0,0.0); 
        (CLK *> O[21])=(0.0,0.0); 
        (CLK *> O[22])=(0.0,0.0); 
        (CLK *> O[23])=(0.0,0.0); 
        (CLK *> O[24])=(0.0,0.0); 
        (CLK *> O[25])=(0.0,0.0); 
        (CLK *> O[26])=(0.0,0.0); 
        (CLK *> O[27])=(0.0,0.0); 
        (CLK *> O[28])=(0.0,0.0); 
        (CLK *> O[29])=(0.0,0.0); 
        (CLK *> O[30])=(0.0,0.0); 
        (CLK *> O[31])=(0.0,0.0); 
      (CLK *> O)=(0.0,0.0);
      (CLK *> ACCUMCO)=(0.0,0.0);
        (ACCUMCI *> O[0])=(0.0,0.0); 
        (ACCUMCI *> O[1])=(0.0,0.0); 
        (ACCUMCI *> O[2])=(0.0,0.0); 
        (ACCUMCI *> O[3])=(0.0,0.0); 
        (ACCUMCI *> O[4])=(0.0,0.0); 
        (ACCUMCI *> O[5])=(0.0,0.0); 
        (ACCUMCI *> O[6])=(0.0,0.0); 
        (ACCUMCI *> O[7])=(0.0,0.0); 
        (ACCUMCI *> O[8])=(0.0,0.0); 
        (ACCUMCI *> O[9])=(0.0,0.0); 
        (ACCUMCI *> O[10])=(0.0,0.0); 
        (ACCUMCI *> O[11])=(0.0,0.0); 
        (ACCUMCI *> O[12])=(0.0,0.0); 
        (ACCUMCI *> O[13])=(0.0,0.0); 
        (ACCUMCI *> O[14])=(0.0,0.0); 
        (ACCUMCI *> O[15])=(0.0,0.0); 
        (ACCUMCI *> O[16])=(0.0,0.0); 
        (ACCUMCI *> O[17])=(0.0,0.0); 
        (ACCUMCI *> O[18])=(0.0,0.0); 
        (ACCUMCI *> O[19])=(0.0,0.0); 
        (ACCUMCI *> O[20])=(0.0,0.0); 
        (ACCUMCI *> O[21])=(0.0,0.0); 
        (ACCUMCI *> O[22])=(0.0,0.0); 
        (ACCUMCI *> O[23])=(0.0,0.0); 
        (ACCUMCI *> O[24])=(0.0,0.0); 
        (ACCUMCI *> O[25])=(0.0,0.0); 
        (ACCUMCI *> O[26])=(0.0,0.0); 
        (ACCUMCI *> O[27])=(0.0,0.0); 
        (ACCUMCI *> O[28])=(0.0,0.0); 
        (ACCUMCI *> O[29])=(0.0,0.0); 
        (ACCUMCI *> O[30])=(0.0,0.0); 
        (ACCUMCI *> O[31])=(0.0,0.0); 
        (ACCUMCI *> O[0])=(0.0,0.0); 
        (ACCUMCI *> O[1])=(0.0,0.0); 
        (ACCUMCI *> O[2])=(0.0,0.0); 
        (ACCUMCI *> O[3])=(0.0,0.0); 
        (ACCUMCI *> O[4])=(0.0,0.0); 
        (ACCUMCI *> O[5])=(0.0,0.0); 
        (ACCUMCI *> O[6])=(0.0,0.0); 
        (ACCUMCI *> O[7])=(0.0,0.0); 
        (ACCUMCI *> O[8])=(0.0,0.0); 
        (ACCUMCI *> O[9])=(0.0,0.0); 
        (ACCUMCI *> O[10])=(0.0,0.0); 
        (ACCUMCI *> O[11])=(0.0,0.0); 
        (ACCUMCI *> O[12])=(0.0,0.0); 
        (ACCUMCI *> O[13])=(0.0,0.0); 
        (ACCUMCI *> O[14])=(0.0,0.0); 
        (ACCUMCI *> O[15])=(0.0,0.0); 
        (ACCUMCI *> O[16])=(0.0,0.0); 
        (ACCUMCI *> O[17])=(0.0,0.0); 
        (ACCUMCI *> O[18])=(0.0,0.0); 
        (ACCUMCI *> O[19])=(0.0,0.0); 
        (ACCUMCI *> O[20])=(0.0,0.0); 
        (ACCUMCI *> O[21])=(0.0,0.0); 
        (ACCUMCI *> O[22])=(0.0,0.0); 
        (ACCUMCI *> O[23])=(0.0,0.0); 
        (ACCUMCI *> O[24])=(0.0,0.0); 
        (ACCUMCI *> O[25])=(0.0,0.0); 
        (ACCUMCI *> O[26])=(0.0,0.0); 
        (ACCUMCI *> O[27])=(0.0,0.0); 
        (ACCUMCI *> O[28])=(0.0,0.0); 
        (ACCUMCI *> O[29])=(0.0,0.0); 
        (ACCUMCI *> O[30])=(0.0,0.0); 
        (ACCUMCI *> O[31])=(0.0,0.0); 
      (ACCUMCI *> CO)=(0.0,0.0);
      (ACCUMCI *> ACCUMCO)=(0.0,0.0);
        (CI *> O[0])=(0.0,0.0); 
        (CI *> O[1])=(0.0,0.0); 
        (CI *> O[2])=(0.0,0.0); 
        (CI *> O[3])=(0.0,0.0); 
        (CI *> O[4])=(0.0,0.0); 
        (CI *> O[5])=(0.0,0.0); 
        (CI *> O[6])=(0.0,0.0); 
        (CI *> O[7])=(0.0,0.0); 
        (CI *> O[8])=(0.0,0.0); 
        (CI *> O[9])=(0.0,0.0); 
        (CI *> O[10])=(0.0,0.0); 
        (CI *> O[11])=(0.0,0.0); 
        (CI *> O[12])=(0.0,0.0); 
        (CI *> O[13])=(0.0,0.0); 
        (CI *> O[14])=(0.0,0.0); 
        (CI *> O[15])=(0.0,0.0); 
        (CI *> O[16])=(0.0,0.0); 
        (CI *> O[17])=(0.0,0.0); 
        (CI *> O[18])=(0.0,0.0); 
        (CI *> O[19])=(0.0,0.0); 
        (CI *> O[20])=(0.0,0.0); 
        (CI *> O[21])=(0.0,0.0); 
        (CI *> O[22])=(0.0,0.0); 
        (CI *> O[23])=(0.0,0.0); 
        (CI *> O[24])=(0.0,0.0); 
        (CI *> O[25])=(0.0,0.0); 
        (CI *> O[26])=(0.0,0.0); 
        (CI *> O[27])=(0.0,0.0); 
        (CI *> O[28])=(0.0,0.0); 
        (CI *> O[29])=(0.0,0.0); 
        (CI *> O[30])=(0.0,0.0); 
        (CI *> O[31])=(0.0,0.0); 
      (CI *> CO)=(0.0,0.0);
      (CI *> ACCUMCO)=(0.0,0.0);
      (CLK *> SIGNEXTOUT)=(0.0,0.0);
        (A[0] *> CO)=(0.0,0.0); 
        (A[1] *> CO)=(0.0,0.0); 
        (A[2] *> CO)=(0.0,0.0); 
        (A[3] *> CO)=(0.0,0.0); 
        (A[4] *> CO)=(0.0,0.0); 
        (A[5] *> CO)=(0.0,0.0); 
        (A[6] *> CO)=(0.0,0.0); 
        (A[7] *> CO)=(0.0,0.0); 
        (A[8] *> CO)=(0.0,0.0); 
        (A[9] *> CO)=(0.0,0.0); 
        (A[10] *> CO)=(0.0,0.0); 
        (A[11] *> CO)=(0.0,0.0); 
        (A[12] *> CO)=(0.0,0.0); 
        (A[13] *> CO)=(0.0,0.0); 
        (A[14] *> CO)=(0.0,0.0); 
        (A[15] *> CO)=(0.0,0.0); 
        (A[0] *> ACCUMCO)=(0.0,0.0); 
        (A[1] *> ACCUMCO)=(0.0,0.0); 
        (A[2] *> ACCUMCO)=(0.0,0.0); 
        (A[3] *> ACCUMCO)=(0.0,0.0); 
        (A[4] *> ACCUMCO)=(0.0,0.0); 
        (A[5] *> ACCUMCO)=(0.0,0.0); 
        (A[6] *> ACCUMCO)=(0.0,0.0); 
        (A[7] *> ACCUMCO)=(0.0,0.0); 
        (A[8] *> ACCUMCO)=(0.0,0.0); 
        (A[9] *> ACCUMCO)=(0.0,0.0); 
        (A[10] *> ACCUMCO)=(0.0,0.0); 
        (A[11] *> ACCUMCO)=(0.0,0.0); 
        (A[12] *> ACCUMCO)=(0.0,0.0); 
        (A[13] *> ACCUMCO)=(0.0,0.0); 
        (A[14] *> ACCUMCO)=(0.0,0.0); 
        (A[15] *> ACCUMCO)=(0.0,0.0); 
        (A[0] *> SIGNEXTOUT)=(0.0,0.0); 
        (A[1] *> SIGNEXTOUT)=(0.0,0.0); 
        (A[2] *> SIGNEXTOUT)=(0.0,0.0); 
        (A[3] *> SIGNEXTOUT)=(0.0,0.0); 
        (A[4] *> SIGNEXTOUT)=(0.0,0.0); 
        (A[5] *> SIGNEXTOUT)=(0.0,0.0); 
        (A[6] *> SIGNEXTOUT)=(0.0,0.0); 
        (A[7] *> SIGNEXTOUT)=(0.0,0.0); 
        (A[8] *> SIGNEXTOUT)=(0.0,0.0); 
        (A[9] *> SIGNEXTOUT)=(0.0,0.0); 
        (A[10] *> SIGNEXTOUT)=(0.0,0.0); 
        (A[11] *> SIGNEXTOUT)=(0.0,0.0); 
        (A[12] *> SIGNEXTOUT)=(0.0,0.0); 
        (A[13] *> SIGNEXTOUT)=(0.0,0.0); 
        (A[14] *> SIGNEXTOUT)=(0.0,0.0); 
        (A[15] *> SIGNEXTOUT)=(0.0,0.0); 
        (D[0] *> CO)=(0.0,0.0); 
        (D[1] *> CO)=(0.0,0.0); 
        (D[2] *> CO)=(0.0,0.0); 
        (D[3] *> CO)=(0.0,0.0); 
        (D[4] *> CO)=(0.0,0.0); 
        (D[5] *> CO)=(0.0,0.0); 
        (D[6] *> CO)=(0.0,0.0); 
        (D[7] *> CO)=(0.0,0.0); 
        (D[8] *> CO)=(0.0,0.0); 
        (D[9] *> CO)=(0.0,0.0); 
        (D[10] *> CO)=(0.0,0.0); 
        (D[11] *> CO)=(0.0,0.0); 
        (D[12] *> CO)=(0.0,0.0); 
        (D[13] *> CO)=(0.0,0.0); 
        (D[14] *> CO)=(0.0,0.0); 
        (D[15] *> CO)=(0.0,0.0); 
        (D[0] *> ACCUMCO)=(0.0,0.0); 
        (D[1] *> ACCUMCO)=(0.0,0.0); 
        (D[2] *> ACCUMCO)=(0.0,0.0); 
        (D[3] *> ACCUMCO)=(0.0,0.0); 
        (D[4] *> ACCUMCO)=(0.0,0.0); 
        (D[5] *> ACCUMCO)=(0.0,0.0); 
        (D[6] *> ACCUMCO)=(0.0,0.0); 
        (D[7] *> ACCUMCO)=(0.0,0.0); 
        (D[8] *> ACCUMCO)=(0.0,0.0); 
        (D[9] *> ACCUMCO)=(0.0,0.0); 
        (D[10] *> ACCUMCO)=(0.0,0.0); 
        (D[11] *> ACCUMCO)=(0.0,0.0); 
        (D[12] *> ACCUMCO)=(0.0,0.0); 
        (D[13] *> ACCUMCO)=(0.0,0.0); 
        (D[14] *> ACCUMCO)=(0.0,0.0); 
        (D[15] *> ACCUMCO)=(0.0,0.0); 
        (D[0] *> SIGNEXTOUT)=(0.0,0.0); 
        (D[1] *> SIGNEXTOUT)=(0.0,0.0); 
        (D[2] *> SIGNEXTOUT)=(0.0,0.0); 
        (D[3] *> SIGNEXTOUT)=(0.0,0.0); 
        (D[4] *> SIGNEXTOUT)=(0.0,0.0); 
        (D[5] *> SIGNEXTOUT)=(0.0,0.0); 
        (D[6] *> SIGNEXTOUT)=(0.0,0.0); 
        (D[7] *> SIGNEXTOUT)=(0.0,0.0); 
        (D[8] *> SIGNEXTOUT)=(0.0,0.0); 
        (D[9] *> SIGNEXTOUT)=(0.0,0.0); 
        (D[10] *> SIGNEXTOUT)=(0.0,0.0); 
        (D[11] *> SIGNEXTOUT)=(0.0,0.0); 
        (D[12] *> SIGNEXTOUT)=(0.0,0.0); 
        (D[13] *> SIGNEXTOUT)=(0.0,0.0); 
        (D[14] *> SIGNEXTOUT)=(0.0,0.0); 
        (D[15] *> SIGNEXTOUT)=(0.0,0.0); 
        (C[0] *> CO)=(0.0,0.0); 
        (C[1] *> CO)=(0.0,0.0); 
        (C[2] *> CO)=(0.0,0.0); 
        (C[3] *> CO)=(0.0,0.0); 
        (C[4] *> CO)=(0.0,0.0); 
        (C[5] *> CO)=(0.0,0.0); 
        (C[6] *> CO)=(0.0,0.0); 
        (C[7] *> CO)=(0.0,0.0); 
        (C[8] *> CO)=(0.0,0.0); 
        (C[9] *> CO)=(0.0,0.0); 
        (C[10] *> CO)=(0.0,0.0); 
        (C[11] *> CO)=(0.0,0.0); 
        (C[12] *> CO)=(0.0,0.0); 
        (C[13] *> CO)=(0.0,0.0); 
        (C[14] *> CO)=(0.0,0.0); 
        (C[15] *> CO)=(0.0,0.0); 
        (C[0] *> ACCUMCO)=(0.0,0.0); 
        (C[1] *> ACCUMCO)=(0.0,0.0); 
        (C[2] *> ACCUMCO)=(0.0,0.0); 
        (C[3] *> ACCUMCO)=(0.0,0.0); 
        (C[4] *> ACCUMCO)=(0.0,0.0); 
        (C[5] *> ACCUMCO)=(0.0,0.0); 
        (C[6] *> ACCUMCO)=(0.0,0.0); 
        (C[7] *> ACCUMCO)=(0.0,0.0); 
        (C[8] *> ACCUMCO)=(0.0,0.0); 
        (C[9] *> ACCUMCO)=(0.0,0.0); 
        (C[10] *> ACCUMCO)=(0.0,0.0); 
        (C[11] *> ACCUMCO)=(0.0,0.0); 
        (C[12] *> ACCUMCO)=(0.0,0.0); 
        (C[13] *> ACCUMCO)=(0.0,0.0); 
        (C[14] *> ACCUMCO)=(0.0,0.0); 
        (C[15] *> ACCUMCO)=(0.0,0.0); 
        (C[0] *> SIGNEXTOUT)=(0.0,0.0); 
        (C[1] *> SIGNEXTOUT)=(0.0,0.0); 
        (C[2] *> SIGNEXTOUT)=(0.0,0.0); 
        (C[3] *> SIGNEXTOUT)=(0.0,0.0); 
        (C[4] *> SIGNEXTOUT)=(0.0,0.0); 
        (C[5] *> SIGNEXTOUT)=(0.0,0.0); 
        (C[6] *> SIGNEXTOUT)=(0.0,0.0); 
        (C[7] *> SIGNEXTOUT)=(0.0,0.0); 
        (C[8] *> SIGNEXTOUT)=(0.0,0.0); 
        (C[9] *> SIGNEXTOUT)=(0.0,0.0); 
        (C[10] *> SIGNEXTOUT)=(0.0,0.0); 
        (C[11] *> SIGNEXTOUT)=(0.0,0.0); 
        (C[12] *> SIGNEXTOUT)=(0.0,0.0); 
        (C[13] *> SIGNEXTOUT)=(0.0,0.0); 
        (C[14] *> SIGNEXTOUT)=(0.0,0.0); 
        (C[15] *> SIGNEXTOUT)=(0.0,0.0); 
        (B[0] *> CO)=(0.0,0.0); 
        (B[1] *> CO)=(0.0,0.0); 
        (B[2] *> CO)=(0.0,0.0); 
        (B[3] *> CO)=(0.0,0.0); 
        (B[4] *> CO)=(0.0,0.0); 
        (B[5] *> CO)=(0.0,0.0); 
        (B[6] *> CO)=(0.0,0.0); 
        (B[7] *> CO)=(0.0,0.0); 
        (B[8] *> CO)=(0.0,0.0); 
        (B[9] *> CO)=(0.0,0.0); 
        (B[10] *> CO)=(0.0,0.0); 
        (B[11] *> CO)=(0.0,0.0); 
        (B[12] *> CO)=(0.0,0.0); 
        (B[13] *> CO)=(0.0,0.0); 
        (B[14] *> CO)=(0.0,0.0); 
        (B[15] *> CO)=(0.0,0.0); 
        (B[0] *> ACCUMCO)=(0.0,0.0); 
        (B[1] *> ACCUMCO)=(0.0,0.0); 
        (B[2] *> ACCUMCO)=(0.0,0.0); 
        (B[3] *> ACCUMCO)=(0.0,0.0); 
        (B[4] *> ACCUMCO)=(0.0,0.0); 
        (B[5] *> ACCUMCO)=(0.0,0.0); 
        (B[6] *> ACCUMCO)=(0.0,0.0); 
        (B[7] *> ACCUMCO)=(0.0,0.0); 
        (B[8] *> ACCUMCO)=(0.0,0.0); 
        (B[9] *> ACCUMCO)=(0.0,0.0); 
        (B[10] *> ACCUMCO)=(0.0,0.0); 
        (B[11] *> ACCUMCO)=(0.0,0.0); 
        (B[12] *> ACCUMCO)=(0.0,0.0); 
        (B[13] *> ACCUMCO)=(0.0,0.0); 
        (B[14] *> ACCUMCO)=(0.0,0.0); 
        (B[15] *> ACCUMCO)=(0.0,0.0); 
        (B[0] *> SIGNEXTOUT)=(0.0,0.0); 
        (B[1] *> SIGNEXTOUT)=(0.0,0.0); 
        (B[2] *> SIGNEXTOUT)=(0.0,0.0); 
        (B[3] *> SIGNEXTOUT)=(0.0,0.0); 
        (B[4] *> SIGNEXTOUT)=(0.0,0.0); 
        (B[5] *> SIGNEXTOUT)=(0.0,0.0); 
        (B[6] *> SIGNEXTOUT)=(0.0,0.0); 
        (B[7] *> SIGNEXTOUT)=(0.0,0.0); 
        (B[8] *> SIGNEXTOUT)=(0.0,0.0); 
        (B[9] *> SIGNEXTOUT)=(0.0,0.0); 
        (B[10] *> SIGNEXTOUT)=(0.0,0.0); 
        (B[11] *> SIGNEXTOUT)=(0.0,0.0); 
        (B[12] *> SIGNEXTOUT)=(0.0,0.0); 
        (B[13] *> SIGNEXTOUT)=(0.0,0.0); 
        (B[14] *> SIGNEXTOUT)=(0.0,0.0); 
        (B[15] *> SIGNEXTOUT)=(0.0,0.0); 
		(CLK *> CO)=(0.0,0.0); 
	 
		  $recovery( posedge IRSTTOP,posedge CLK , 1.0);
		  $recovery( negedge IRSTTOP, posedge CLK ,1.0);   
		  $removal( posedge IRSTTOP, posedge CLK ,1.0);
		  $removal( negedge IRSTTOP, posedge CLK ,1.0);
		  $recovery(posedge IRSTBOT , posedge CLK ,1.0);
		  $recovery(negedge IRSTBOT , posedge CLK ,1.0);	 
		  $removal(posedge IRSTBOT , posedge CLK ,1.0);
		  $removal(negedge IRSTBOT , posedge CLK ,1.0);
		  $recovery( posedge ORSTTOP, posedge CLK ,1.0);
		  $recovery( negedge ORSTTOP, posedge CLK ,1.0);
		  $removal( posedge ORSTTOP, posedge CLK ,1.0);
		  $removal( negedge ORSTTOP, posedge CLK ,1.0);
		  $recovery(posedge ORSTBOT , posedge CLK ,1.0);
		  $recovery(negedge ORSTBOT , posedge CLK ,1.0);	   
		  $removal(posedge ORSTBOT , posedge CLK ,1.0);
		  $removal(negedge ORSTBOT , posedge CLK ,1.0);
		  $width (posedge CLK, 1.0 ); 
		  $period (posedge CLK, 1.0 ); 

		  $setuphold( posedge CLK,posedge A[0],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge A[0],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge A[1],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge A[1],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge A[2],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge A[2],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge A[3],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge A[3],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge A[4],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge A[4],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge A[5],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge A[5],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge A[6],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge A[6],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge A[7],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge A[7],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge A[8],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge A[8],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge A[9],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge A[9],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge A[10],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge A[10],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge A[11],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge A[11],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge A[12],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge A[12],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge A[13],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge A[13],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge A[14],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge A[14],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge A[15],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge A[15],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge B[0],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge B[0],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge B[1],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge B[1],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge B[2],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge B[2],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge B[3],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge B[3],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge B[4],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge B[4],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge B[5],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge B[5],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge B[6],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge B[6],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge B[7],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge B[7],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge B[8],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge B[8],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge B[9],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge B[9],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge B[10],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge B[10],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge B[11],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge B[11],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge B[12],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge B[12],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge B[13],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge B[13],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge B[14],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge B[14],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge B[15],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge B[15],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge C[0],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge C[0],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge C[1],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge C[1],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge C[2],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge C[2],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge C[3],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge C[3],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge C[4],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge C[4],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge C[5],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge C[5],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge C[6],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge C[6],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge C[7],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge C[7],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge C[8],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge C[8],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge C[9],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge C[9],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge C[10],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge C[10],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge C[11],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge C[11],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge C[12],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge C[12],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge C[13],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge C[13],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge C[14],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge C[14],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge C[15],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge C[15],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge D[0],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge D[0],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge D[1],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge D[1],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge D[2],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge D[2],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge D[3],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge D[3],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge D[4],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge D[4],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge D[5],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge D[5],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge D[6],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge D[6],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge D[7],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge D[7],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge D[8],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge D[8],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge D[9],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge D[9],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge D[10],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge D[10],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge D[11],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge D[11],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge D[12],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge D[12],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge D[13],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge D[13],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge D[14],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge D[14],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge D[15],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge D[15],1.0, 1.0, NOTIFIER);
		  
		  
		  
		
		   $setuphold(posedge CLK, posedge AHOLD, 1.0, 1.0, NOTIFIER);
		   $setuphold(posedge CLK, posedge BHOLD, 1.0, 1.0, NOTIFIER);
		   $setuphold(posedge CLK, posedge CHOLD, 1.0, 1.0, NOTIFIER);
		   $setuphold(posedge CLK, posedge DHOLD, 1.0, 1.0, NOTIFIER);
		   $setuphold(posedge CLK, posedge ADDSUBTOP, 1.0, 1.0, NOTIFIER);
		   $setuphold(posedge CLK, posedge OHOLDTOP, 1.0, 1.0, NOTIFIER);
		   $setuphold(posedge CLK, posedge ADDSUBBOT, 1.0, 1.0, NOTIFIER);
		   $setuphold(posedge CLK, posedge OHOLDBOT, 1.0, 1.0, NOTIFIER);
		   $setuphold(posedge CLK, posedge OLOADTOP, 1.0, 1.0, NOTIFIER);
		   $setuphold(posedge CLK, posedge OLOADBOT, 1.0, 1.0, NOTIFIER);
		   $setuphold(posedge CLK, posedge CI, 1.0, 1.0, NOTIFIER);
		   $setuphold(posedge CLK, posedge ACCUMCI, 1.0, 1.0, NOTIFIER);	 
		   
		  
		   $setuphold(posedge CLK, negedge AHOLD, 1.0, 1.0, NOTIFIER);
		   $setuphold(posedge CLK, negedge BHOLD, 1.0, 1.0, NOTIFIER);
		   $setuphold(posedge CLK, negedge CHOLD, 1.0, 1.0, NOTIFIER);
		   $setuphold(posedge CLK, negedge DHOLD, 1.0, 1.0, NOTIFIER);
		   $setuphold(posedge CLK, negedge ADDSUBTOP, 1.0, 1.0, NOTIFIER);
		   $setuphold(posedge CLK, negedge OHOLDTOP, 1.0, 1.0, NOTIFIER);
		   $setuphold(posedge CLK, negedge ADDSUBBOT, 1.0, 1.0, NOTIFIER);
		   $setuphold(posedge CLK, negedge OHOLDBOT, 1.0, 1.0, NOTIFIER);
		   $setuphold(posedge CLK, negedge OLOADTOP, 1.0, 1.0, NOTIFIER);
		   $setuphold(posedge CLK, negedge OLOADBOT, 1.0, 1.0, NOTIFIER);
		   $setuphold(posedge CLK, negedge CI, 1.0, 1.0, NOTIFIER);
		   $setuphold(posedge CLK, negedge ACCUMCI, 1.0, 1.0, NOTIFIER);
 
		 
		 
		 
		 endspecify
`endif		   
		

endmodule

//////////////////////////////////////////////////////////////////////////////////
// mac16_physical
//////////////////////////////////////////////////////////////////////////////////

`timescale 1ns / 1ps

module mac16_physical  (
	 CLK ,
	 IHRST,
	 ILRST,
	 OHRST,
	 OLRST,
	 
	 A ,
	 B ,
	 C ,
	 D ,
	 
	 CBIT,
	 
	 AHLD,
	 BHLD,
	 CHLD,
	 DHLD,
	 OHHLD,
	 OLHLD,

 
	 OHADS,
	 OLADS,
	 OHLDA,
	 OLLDA,
	 
	 CICAS,
	 CI,
	 SIGNEXTIN,
	 SIGNEXTOUT,

	 COCAS,
	 CO,
	 O
    );

	 input CLK ;
	 input IHRST;
	 input ILRST;
	 input OHRST;
	 input OLRST;
	 
	 input [15:0] A ;
	 input [15:0] B ;
	 input [15:0] C ;
	 input [15:0] D ;
	 
	 input [24:0] CBIT;
	 
	 input AHLD;
	 input BHLD;
	 input CHLD;
	 input DHLD;
	 input OHHLD;
	 input OLHLD;

 
	 input OHADS;
	 input OLADS;
	 input OHLDA;
	 input OLLDA;
	 
	 input CICAS;
	 input CI;
	 input SIGNEXTIN;
	 output SIGNEXTOUT;
	 
	 output COCAS;
	 output CO;
	 output [31:0] O;
	
	
wire AENA, BENA, CENA, DENA, OHENA, OLENA;
assign AENA = ~AHLD;
assign BENA = ~BHLD;
assign CENA = ~CHLD;
assign DENA = ~DHLD;

assign OHENA = ~OHHLD;
assign OLENA = ~OLHLD;


wire ASEL, BSEL, CSEL, DSEL, FSEL, JKSEL, GSEL, HSEL;
wire OHADDA_SEL, OLADDA_SEL, MPY_8X8_MODE, ASGND, BSGND;
wire [1:0] OHOMUX_SEL, OLOMUX_SEL, OHADDB_SEL, OLADDB_SEL, OHCARRYMUX_SEL, OLCARRYMUX_SEL;

assign ASEL = CBIT[1];
assign BSEL = CBIT[2];
assign CSEL = CBIT[0];
assign DSEL = CBIT[3];

assign FSEL = CBIT[4];
assign JKSEL = CBIT[6];
assign GSEL = CBIT[5];
assign HSEL = CBIT[7];

assign OHOMUX_SEL[1:0] = CBIT[9:8];	
assign OLOMUX_SEL[1:0] = CBIT[16:15];	
assign OHADDA_SEL = CBIT[12];
assign OLADDA_SEL = CBIT[19];
assign OHADDB_SEL[1:0] = CBIT[11:10];	
assign OLADDB_SEL[1:0] = CBIT[18:17];	
assign OHCARRYMUX_SEL[1:0] = CBIT[14:13];
assign OLCARRYMUX_SEL[1:0] = CBIT[21:20];
assign MPY_8X8_MODE = CBIT[22];
assign ASGND = CBIT[23];
assign BSGND = CBIT[24];

wire [15:0] REG_A ;
wire [15:0] REG_B ;
wire [15:0] REG_C ;
wire [15:0] REG_D ;

wire [15:0] OH_8X8;
wire [15:0] OL_8X8;
wire [31:0] O_16X16;

wire MAC16_SIGNOUT_L, MAC16_SIGNOUT_H;

assign SIGNEXTOUT = MAC16_SIGNOUT_H;

REG_BYPASS_MUX  A_REG (
	.D(A) ,
	.Q(REG_A) ,
	.ENA(AENA) ,
	.CLK(CLK) ,
	.RST(IHRST) ,
	.SELM(ASEL) 
); 

REG_BYPASS_MUX  B_REG (
	.D(B) ,
	.Q(REG_B) ,
	.ENA(BENA) ,
	.CLK(CLK) ,
	.RST(ILRST) ,
	.SELM(BSEL) 
); 

REG_BYPASS_MUX  C_REG (
	.D(C) ,
	.Q(REG_C) ,
	.ENA(CENA) ,
	.CLK(CLK) ,
	.RST(IHRST) ,
	.SELM(CSEL) 
); 

REG_BYPASS_MUX  D_REG (
	.D(D) ,
	.Q(REG_D) ,
	.ENA(DENA) ,
	.CLK(CLK) ,
	.RST(ILRST) ,
	.SELM(DSEL) 
); 

MULT_ACCUM HI_MAC (
	.DIRECT_INPUT(REG_C),
	.MULT_INPUT(REG_A),
	.MULT_8x8(OH_8X8[15:0]),
	.MULT_16x16(O_16X16[31:16]),
	.ADDSUB(OHADS),
	.CLK(CLK),
	.CICAS(COCAS_L),
	.CI(CO_L),
	.SIGNEXTIN(MAC16_SIGNOUT_L) ,
	.SIGNEXTOUT(MAC16_SIGNOUT_H) ,
	.LDA(OHLDA),
	.RST(OHRST),
	.ENA(OHENA),
	.COCAS(COCAS),
	.CO(CO),
	.O(O[31:16]),
	.OUTMUX_SEL(OHOMUX_SEL[1:0]),
	.ADDER_A_IN_SEL(OHADDA_SEL),
	.ADDER_B_IN_SEL(OHADDB_SEL[1:0]),
	.CARRYMUX_SEL(OHCARRYMUX_SEL[1:0])
    );

MULT_ACCUM LO_MAC (
	.DIRECT_INPUT(REG_D),
	.MULT_INPUT(REG_B),
	.MULT_8x8(OL_8X8[15:0]),
	.MULT_16x16(O_16X16[15:0]),
	.ADDSUB(OLADS),
	.CLK(CLK),
	.CICAS(CICAS),
	.CI(CI),
	.SIGNEXTIN(SIGNEXTIN) ,
	.SIGNEXTOUT(MAC16_SIGNOUT_L) ,
	.LDA(OLLDA),
	.RST(OLRST),
	.ENA(OLENA),
	.COCAS(COCAS_L),
	.CO(CO_L),
	.O(O[15:0]),
	.OUTMUX_SEL(OLOMUX_SEL[1:0]),
	.ADDER_A_IN_SEL(OLADDA_SEL),
	.ADDER_B_IN_SEL(OLADDB_SEL[1:0]),
	.CARRYMUX_SEL(OLCARRYMUX_SEL[1:0])
    );
	 
MPY16X16 MULTIPLER (
	.clk(CLK),
	.IHRST(IHRST),
	.ILRST(ILRST),
	.FSEL(FSEL),
	.GSEL(GSEL),
	.HSEL(HSEL),
	.JKSEL(JKSEL),
	.MPY_8X8_MODE(MPY_8X8_MODE),
	.ASGND(ASGND),
	.BSGND(BSGND),
	.A(REG_A[15:0]),
	.B(REG_B[15:0]),
	.OH_8X8(OH_8X8[15:0]),
	.OL_8X8(OL_8X8[15:0]),
	.O_16X16(O_16X16[31:0])
);

endmodule


//////////////////////////////////////////////////////////////////////////////////
// Module Name:    MPY16X16
//////////////////////////////////////////////////////////////////////////////////

`timescale 1ns / 1ps

//////////////////////////////////////////////////// 
`define  SIGNED_DATA		1'b1
`define  UNSIGNED_DATA		1'b0
////////////////////////////////////////////////////

module booth_encoder(booth_single, booth_double, booth_negtive, multiplier, signed_mpy);
input	[7:0]multiplier;
output	[4:0]booth_single;
output	[4:0]booth_double;
output	[4:0]booth_negtive;
input	signed_mpy;

wire	[10:0]booth_in;
wire	[1:0]sign_ext;
assign sign_ext=(signed_mpy==1'b1)?{2{multiplier[7]}} : 2'b00;

assign booth_in={sign_ext ,multiplier[7:0],1'b0};


assign  booth_negtive[0]=booth_in[2];
assign  booth_negtive[1]=booth_in[4];
assign  booth_negtive[2]=booth_in[6];
assign  booth_negtive[3]=booth_in[8];
assign  booth_negtive[4]=booth_in[10];

assign  booth_single[0]=booth_in[0]^booth_in[1];
assign  booth_single[1]=booth_in[2]^booth_in[3];
assign  booth_single[2]=booth_in[4]^booth_in[5];
assign  booth_single[3]=booth_in[6]^booth_in[7];
assign  booth_single[4]=booth_in[8]^booth_in[9];


assign  booth_double[0]=~(~(booth_in[0] & booth_in[1] & ~booth_in[2]) & ~(~booth_in[0] & ~booth_in[1] & booth_in[2]));
assign  booth_double[1]=~(~(booth_in[2] & booth_in[3] & ~booth_in[4]) & ~(~booth_in[2] & ~booth_in[3] & booth_in[4]));
assign  booth_double[2]=~(~(booth_in[4] & booth_in[5] & ~booth_in[6]) & ~(~booth_in[4] & ~booth_in[5] & booth_in[6]));
assign  booth_double[3]=~(~(booth_in[6] & booth_in[7] & ~booth_in[8]) & ~(~booth_in[6] & ~booth_in[7] & booth_in[8]));
assign  booth_double[4]=~(~(booth_in[8] & booth_in[9] & ~booth_in[10]) & ~(~booth_in[8] & ~booth_in[9] & booth_in[10]));

endmodule // booth_encoder

///////////////////////////////////////////////////////////////////////

`timescale 1ns / 1ps 

module booth_selector(pp_out,booth_single, booth_double, booth_negtive,multiplicand, signed_mpy);
input	[7:0]multiplicand;
input	[4:0]booth_single;
input	[4:0]booth_double;
input	[4:0]booth_negtive;
output	[44:0] pp_out;
integer	j;

reg		[8:0] pp0,pp1,pp2,pp3,pp4;

input	signed_mpy;
wire	sign_ext;
assign sign_ext=(signed_mpy==1'b1)?{multiplicand[7]} : 1'b0;


assign pp_out ={pp4, pp3, pp2, pp1, pp0};

wire	[9:0]bs_in;

assign  bs_in={sign_ext ,multiplicand[7:0],1'b0};


always @(booth_negtive or booth_single or bs_in or booth_double)

begin
	for (j=0; j<=8; j=j+1)
	begin
		pp0[j] = (booth_negtive[0]^ ~(~(booth_single[0] & bs_in[j+1]) & ~(booth_double[0] & bs_in[j])));
		pp1[j] = (booth_negtive[1]^ ~(~(booth_single[1] & bs_in[j+1]) & ~(booth_double[1] & bs_in[j])));
		pp2[j] = (booth_negtive[2]^ ~(~(booth_single[2] & bs_in[j+1]) & ~(booth_double[2] & bs_in[j])));
		pp3[j] = (booth_negtive[3]^ ~(~(booth_single[3] & bs_in[j+1]) & ~(booth_double[3] & bs_in[j])));
		pp4[j] = (booth_negtive[4]^ ~(~(booth_single[4] & bs_in[j+1]) & ~(booth_double[4] & bs_in[j])));
	end

end 

endmodule // booth_selector

///////////////////////////////////////////////////////////////////////
`timescale 1ns / 1ps

module MPY8x8(csa_a,csa_b,multiplicand,multiplier,signed_MPD,signed_MPR);
input	[7:0]multiplicand;
input	[7:0]multiplier;
input	signed_MPD, signed_MPR;

output [15:0] csa_a;
output [15:0] csa_b;

wire	[4:0]booth_single;
wire	[4:0]booth_double;
wire	[4:0]booth_negtive;
wire	[4:0]pp_sign;

wire	[44:0]pp_out;
wire	[8:0] PP0,PP1,PP2,PP3,PP4;

assign {PP4, PP3, PP2, PP1, PP0} = pp_out;

booth_encoder booth_encoder
(
.booth_single(booth_single), 
.booth_double(booth_double), 
.booth_negtive(booth_negtive), 
.multiplier(multiplier),
.signed_mpy(signed_MPR)
);


booth_selector booth_selector
(
.pp_out(pp_out),
.booth_single(booth_single), 
.booth_double(booth_double), 
.booth_negtive(booth_negtive),
.multiplicand(multiplicand),
.signed_mpy(signed_MPD)
);

wire	current_MPD_sign;
assign current_MPD_sign = multiplicand[7] & signed_MPD;
//assign pp_sign[0] = (booth_negtive[0] ^ current_MPD_sign) & (booth_single[0] | booth_double[0] | booth_negtive[0]) | (~booth_single[0] & ~booth_double[0] & booth_negtive[0]);
//assign pp_sign[1] = (booth_negtive[1] ^ current_MPD_sign) & (booth_single[1] | booth_double[1] | booth_negtive[1]) | (~booth_single[1] & ~booth_double[1] & booth_negtive[1]);
//assign pp_sign[2] = (booth_negtive[2] ^ current_MPD_sign) & (booth_single[2] | booth_double[2] | booth_negtive[2]) | (~booth_single[2] & ~booth_double[2] & booth_negtive[2]);
//assign pp_sign[3] = (booth_negtive[3] ^ current_MPD_sign) & (booth_single[3] | booth_double[3] | booth_negtive[3]) | (~booth_single[3] & ~booth_double[3] & booth_negtive[3]);
//assign pp_sign[4] = (booth_negtive[4] ^ current_MPD_sign) & (booth_single[4] | booth_double[4] | booth_negtive[4]) | (~booth_single[4] & ~booth_double[4] & booth_negtive[4]);

integer j;
reg [4:0] booth_single_b, booth_double_b, booth_negtive_b;

always @(booth_single or booth_double or booth_negtive)
begin
	for (j=0; j<=4; j=j+1)
	begin
		booth_single_b[j] = ~booth_single[j];
		booth_double_b[j] = ~booth_double[j];
		booth_negtive_b[j] = ~booth_negtive[j];
	end
end 

assign pp_sign[0] = (booth_negtive[0] ^ current_MPD_sign) & ~(booth_single_b[0] & booth_double_b[0] & booth_negtive_b[0]) | (booth_single_b[0] & booth_double_b[0] & booth_negtive[0]);
assign pp_sign[1] = (booth_negtive[1] ^ current_MPD_sign) & ~(booth_single_b[1] & booth_double_b[1] & booth_negtive_b[1]) | (booth_single_b[1] & booth_double_b[1] & booth_negtive[1]);
assign pp_sign[2] = (booth_negtive[2] ^ current_MPD_sign) & ~(booth_single_b[2] & booth_double_b[2] & booth_negtive_b[2]) | (booth_single_b[2] & booth_double_b[2] & booth_negtive[2]);
assign pp_sign[3] = (booth_negtive[3] ^ current_MPD_sign) & ~(booth_single_b[3] & booth_double_b[3] & booth_negtive_b[3]) | (booth_single_b[3] & booth_double_b[3] & booth_negtive[3]);
assign pp_sign[4] = (booth_negtive[4] ^ current_MPD_sign) & ~(booth_single_b[4] & booth_double_b[4] & booth_negtive_b[4]) | (booth_single_b[4] & booth_double_b[4] & booth_negtive[4]);
// Wallace CSA step#1

wire	FA1_R00C14_C, FA1_R00C14_S;
wire	FA1_R00C13_C, FA1_R00C13_S;
wire	FA1_R00C12_C, FA1_R00C12_S;

wire	FA1_R00C11_C, FA1_R00C11_S;
wire	HA1_R03C11_C, HA1_R03C11_S;

wire	FA1_R00C10_C, FA1_R00C10_S;
wire	HA1_R03C10_C, HA1_R03C10_S;

wire	FA1_R00C09_C, FA1_R00C09_S;
wire	HA1_R03C09_C, HA1_R03C09_S;

wire	FA1_R00C08_C, FA1_R00C08_S;
wire	FA1_R03C08_C, FA1_R03C08_S;

wire	FA1_R00C07_C, FA1_R00C07_S;
wire	FA1_R00C06_C, FA1_R00C06_S;
wire	HA1_R03C06_C, HA1_R03C06_S;

wire	FA1_R00C05_C, FA1_R00C05_S;
wire	FA1_R00C04_C, FA1_R00C04_S;

wire	FA1_R00C02_C, FA1_R00C02_S;


fa FA1_R00C14(.Cout(FA1_R00C14_C), .Sum(FA1_R00C14_S), .A(1'b1), .B(PP3[8]), .C(PP4[6]));

fa FA1_R00C13(.Cout(FA1_R00C13_C), .Sum(FA1_R00C13_S), .A(~pp_sign[2]), .B(PP3[7]), .C(PP4[5]));

fa FA1_R00C12(.Cout(FA1_R00C12_C), .Sum(FA1_R00C12_S), .A(1'b1), .B(PP2[8]), .C(PP3[6]));

fa FA1_R00C11(.Cout(FA1_R00C11_C), .Sum(FA1_R00C11_S), .A(~pp_sign[0]), .B(~pp_sign[1]), .C(PP2[7]));
ha HA1_R03C11(.Cout(HA1_R03C11_C), .Sum(HA1_R03C11_S), .A(PP3[5]), .B(PP4[3]));

fa FA1_R00C10(.Cout(FA1_R00C10_C), .Sum(FA1_R00C10_S), .A(pp_sign[0]), .B(PP1[8]), .C(PP2[6]));
ha HA1_R03C10(.Cout(HA1_R03C10_C), .Sum(HA1_R03C10_S), .A(PP3[4]), .B(PP4[2]));

fa FA1_R00C09(.Cout(FA1_R00C09_C), .Sum(FA1_R00C09_S), .A(pp_sign[0]), .B(PP1[7]), .C(PP2[5]));
ha HA1_R03C09(.Cout(HA1_R03C09_C), .Sum(HA1_R03C09_S), .A(PP3[3]), .B(PP4[1]));

fa FA1_R00C08(.Cout(FA1_R00C08_C), .Sum(FA1_R00C08_S), .A(PP0[8]), .B(PP1[6]), .C(PP2[4]));
fa FA1_R03C08(.Cout(FA1_R03C08_C), .Sum(FA1_R03C08_S), .A(PP3[2]), .B(PP4[0]), .C(booth_negtive[4]));

fa FA1_R00C07(.Cout(FA1_R00C07_C), .Sum(FA1_R00C07_S), .A(PP0[7]), .B(PP1[5]), .C(PP2[3]));
fa FA1_R00C06(.Cout(FA1_R00C06_C), .Sum(FA1_R00C06_S), .A(PP0[6]), .B(PP1[4]), .C(PP2[2]));
ha HA1_R03C06(.Cout(HA1_R03C06_C), .Sum(HA1_R03C06_S), .A(PP3[0]), .B(booth_negtive[3]));

fa FA1_R00C05(.Cout(FA1_R00C05_C), .Sum(FA1_R00C05_S), .A(PP0[5]), .B(PP1[3]), .C(PP2[1]));
fa FA1_R00C04(.Cout(FA1_R00C04_C), .Sum(FA1_R00C04_S), .A(PP0[4]), .B(PP1[2]), .C(PP2[0]));

fa FA1_R00C02(.Cout(FA1_R00C02_C), .Sum(FA1_R00C02_S), .A(PP0[2]), .B(PP1[0]), .C(booth_negtive[1]));

// Wallace CSA step#2

wire	FA2_R00C15_C, FA2_R00C15_S;
wire	HA2_R00C14_C, HA2_R00C14_S;
wire	HA2_R00C13_C, HA2_R00C13_S;

wire	FA2_R00C12_C, FA2_R00C12_S;
wire	FA2_R00C11_C, FA2_R00C11_S;
wire	FA2_R00C10_C, FA2_R00C10_S;
wire	FA2_R00C09_C, FA2_R00C09_S;
wire	FA2_R00C08_C, FA2_R00C08_S;
wire	FA2_R00C07_C, FA2_R00C07_S;
wire	FA2_R00C06_C, FA2_R00C06_S;

wire	FA2_R00C03_C, FA2_R00C03_S;


fa FA2_R00C15(.Cout(FA2_R00C15_C), .Sum(FA2_R00C15_S), .A(~pp_sign[3]), .B(PP4[7]), .C(FA1_R00C14_C));

ha HA2_R00C14(.Cout(HA2_R00C14_C), .Sum(HA2_R00C14_S), .A(FA1_R00C14_S), .B(FA1_R00C13_C));
ha HA2_R00C13(.Cout(HA2_R00C13_C), .Sum(HA2_R00C13_S), .A(FA1_R00C13_S), .B(FA1_R00C12_C));

fa FA2_R00C12(.Cout(FA2_R00C12_C), .Sum(FA2_R00C12_S), .A(FA1_R00C12_S), .B(FA1_R00C11_C), .C(HA1_R03C11_C));
fa FA2_R00C11(.Cout(FA2_R00C11_C), .Sum(FA2_R00C11_S), .A(FA1_R00C11_S), .B(FA1_R00C10_C), .C(HA1_R03C11_S));
fa FA2_R00C10(.Cout(FA2_R00C10_C), .Sum(FA2_R00C10_S), .A(FA1_R00C10_S), .B(FA1_R00C09_C), .C(HA1_R03C10_S));
fa FA2_R00C09(.Cout(FA2_R00C09_C), .Sum(FA2_R00C09_S), .A(FA1_R00C09_S), .B(FA1_R00C08_C), .C(HA1_R03C09_S));
fa FA2_R00C08(.Cout(FA2_R00C08_C), .Sum(FA2_R00C08_S), .A(FA1_R00C08_S), .B(FA1_R00C07_C), .C(FA1_R03C08_S));
fa FA2_R00C07(.Cout(FA2_R00C07_C), .Sum(FA2_R00C07_S), .A(FA1_R00C07_S), .B(FA1_R00C06_C), .C(HA1_R03C06_C));
fa FA2_R00C06(.Cout(FA2_R00C06_C), .Sum(FA2_R00C06_S), .A(FA1_R00C06_S), .B(FA1_R00C05_C), .C(HA1_R03C06_S));

fa FA2_R00C03(.Cout(FA2_R00C03_C), .Sum(FA2_R00C03_S), .A(PP0[3]), .B(PP1[1]), .C(FA1_R00C02_C));

// Wallace CSA step#3
wire	HA3_R00C15_C, HA3_R00C15_S;
wire	HA3_R00C14_C, HA3_R00C14_S;
wire	HA3_R00C13_C, HA3_R00C13_S;
wire	FA3_R00C12_C, FA3_R00C12_S;
wire	FA3_R00C11_C, FA3_R00C11_S;
wire	FA3_R00C10_C, FA3_R00C10_S;
wire	FA3_R00C09_C, FA3_R00C09_S;

wire	HA3_R00C08_C, HA3_R00C08_S;
wire	FA3_R00C07_C, FA3_R00C07_S;

wire	HA3_R00C05_C, HA3_R00C05_S;
wire	FA3_R00C04_C, FA3_R00C04_S;


ha HA3_R00C15(.Cout(HA3_R00C15_C), .Sum(HA3_R00C15_S), .A(FA2_R00C15_S), .B(HA2_R00C14_C));
ha HA3_R00C14(.Cout(HA3_R00C14_C), .Sum(HA3_R00C14_S), .A(HA2_R00C14_S), .B(HA2_R00C13_C));
ha HA3_R00C13(.Cout(HA3_R00C13_C), .Sum(HA3_R00C13_S), .A(HA2_R00C13_S), .B(FA2_R00C12_C));
fa FA3_R00C12(.Cout(FA3_R00C12_C), .Sum(FA3_R00C12_S), .A(FA2_R00C12_S), .B(FA2_R00C11_C), .C(PP4[4]));
fa FA3_R00C11(.Cout(FA3_R00C11_C), .Sum(FA3_R00C11_S), .A(FA2_R00C11_S), .B(FA2_R00C10_C), .C(HA1_R03C10_C));
fa FA3_R00C10(.Cout(FA3_R00C10_C), .Sum(FA3_R00C10_S), .A(FA2_R00C10_S), .B(FA2_R00C09_C), .C(HA1_R03C09_C));
fa FA3_R00C09(.Cout(FA3_R00C09_C), .Sum(FA3_R00C09_S), .A(FA2_R00C09_S), .B(FA2_R00C08_C), .C(FA1_R03C08_C));

ha HA3_R00C08(.Cout(HA3_R00C08_C), .Sum(HA3_R00C08_S), .A(FA2_R00C08_S), .B(FA2_R00C07_C));
fa FA3_R00C07(.Cout(FA3_R00C07_C), .Sum(FA3_R00C07_S), .A(FA2_R00C07_S), .B(FA2_R00C06_C), .C(PP3[1]));

ha HA3_R00C05(.Cout(HA3_R00C05_C), .Sum(HA3_R00C05_S), .A(FA1_R00C05_S), .B(FA1_R00C04_C));
fa FA3_R00C04(.Cout(FA3_R00C04_C), .Sum(FA3_R00C04_S), .A(FA1_R00C04_S), .B(booth_negtive[2]), .C(FA2_R00C03_C));


assign csa_a[0] = PP0[0];
assign csa_b[0] = booth_negtive[0];
assign csa_a[1] = PP0[1];
assign csa_b[1] = 1'b0;
assign csa_a[2] = FA1_R00C02_S;
assign csa_b[2] = 1'b0;
assign csa_a[3] = FA2_R00C03_S;
assign csa_b[3] = 1'b0;

assign csa_a[4] = FA3_R00C04_S;
assign csa_b[4] = 1'b0;

assign csa_a[5] = HA3_R00C05_S;
assign csa_b[5] = FA3_R00C04_C;
assign csa_a[6] = FA2_R00C06_S;
assign csa_b[6] = HA3_R00C05_C;
assign csa_a[7] = FA3_R00C07_S;
assign csa_b[7] = 1'b0;
assign csa_a[8] = HA3_R00C08_S;
assign csa_b[8] = FA3_R00C07_C;
assign csa_a[9] = FA3_R00C09_S;
assign csa_b[9] = HA3_R00C08_C;
assign csa_a[10] = FA3_R00C10_S;
assign csa_b[10] = FA3_R00C09_C;
assign csa_a[11] = FA3_R00C11_S;
assign csa_b[11] = FA3_R00C10_C;
assign csa_a[12] = FA3_R00C12_S;
assign csa_b[12] = FA3_R00C11_C;
assign csa_a[13] = HA3_R00C13_S;
assign csa_b[13] = FA3_R00C12_C;
assign csa_a[14] = HA3_R00C14_S;
assign csa_b[14] = HA3_R00C13_C;
assign csa_a[15] = HA3_R00C15_S;
assign csa_b[15] = HA3_R00C14_C;

endmodule // MPY8x8

///////////////////////////////////////////////////////////////////////
`timescale 1ns / 1ps
module MPY16X16(
clk,

IHRST,
ILRST,

FSEL,
GSEL,
HSEL,
JKSEL,
MPY_8X8_MODE,

ASGND,
BSGND,

A,
B,

OH_8X8,
OL_8X8,
O_16X16
);

input clk;

input IHRST;
input ILRST;

input FSEL;
input GSEL;
input HSEL;
input JKSEL;
input MPY_8X8_MODE;

input ASGND;
input BSGND;

input	[15:0]A;
input	[15:0]B;

output [15:0] OH_8X8;
output [15:0] OL_8X8;
output [31:0] O_16X16;


reg 	[31:0]csa_rega, csa_regb;
wire	[152:0]pp_out;

wire	[7:0] MPYG_mpd, MPYG_mpr;
wire	[7:0] MPYJ_mpd, MPYJ_mpr;
wire	[7:0] MPYF_mpd, MPYF_mpr;
wire	[7:0] MPYK_mpd, MPYK_mpr;

wire	MPYG_MPD_sign, MPYG_MPR_sign;
wire	MPYJ_MPD_sign, MPYJ_MPR_sign;
wire	MPYF_MPD_sign, MPYF_MPR_sign;
wire	MPYK_MPD_sign, MPYK_MPR_sign;

assign MPYG_mpd = A[7:0];
assign MPYG_mpr = B[7:0];
assign MPYG_MPD_sign = MPY_8X8_MODE ? ASGND : `UNSIGNED_DATA;
assign MPYG_MPR_sign = MPY_8X8_MODE ? BSGND : `UNSIGNED_DATA;

assign MPYJ_mpd = A[7:0];
assign MPYJ_mpr = B[15:8];
assign MPYJ_MPD_sign = `UNSIGNED_DATA;
assign MPYJ_MPR_sign = BSGND;

assign MPYF_mpd = A[15:8];
assign MPYF_mpr = B[15:8];
assign MPYF_MPD_sign = ASGND;
assign MPYF_MPR_sign = BSGND;

assign MPYK_mpd = A[15:8];
assign MPYK_mpr = B[7:0];
assign MPYK_MPD_sign = ASGND;
assign MPYK_MPR_sign = `UNSIGNED_DATA;

wire	[15:0] MPYG_csa_a, MPYG_csa_b;
wire	[15:0] MPYJ_csa_a, MPYJ_csa_b;
wire	[15:0] MPYF_csa_a, MPYF_csa_b;
wire	[15:0] MPYK_csa_a, MPYK_csa_b;

wire	[15:0] MPYG_o, MPYG_out;
wire	[15:0] MPYJ_o, MPYJ_out;
wire	[15:0] MPYF_o, MPYF_out;
wire	[15:0] MPYK_o, MPYK_out;
reg		[15:0] MPYG_oreg, MPYJ_oreg;
reg		[15:0] MPYF_oreg, MPYK_oreg;

wire	MPYJ_out_sign, MPYK_out_sign;
wire	MPYJK_g, MPYJK_p;

assign MPYJ_out_sign = BSGND ? MPYJ_out[15] : `UNSIGNED_DATA;
assign MPYK_out_sign = ASGND ? MPYK_out[15] : `UNSIGNED_DATA;

assign MPYJK_g = MPYJ_out_sign & MPYK_out_sign;
assign MPYJK_p = MPYJ_out_sign ^ MPYK_out_sign;


MPY8x8 MPY_G(.csa_a(MPYG_csa_a),.csa_b(MPYG_csa_b),.multiplicand(MPYG_mpd),.multiplier(MPYG_mpr),.signed_MPD(MPYG_MPD_sign),.signed_MPR(MPYG_MPR_sign));
MPY8x8 MPY_J(.csa_a(MPYJ_csa_a),.csa_b(MPYJ_csa_b),.multiplicand(MPYJ_mpd),.multiplier(MPYJ_mpr),.signed_MPD(MPYJ_MPD_sign),.signed_MPR(MPYJ_MPR_sign));
MPY8x8 MPY_F(.csa_a(MPYF_csa_a),.csa_b(MPYF_csa_b),.multiplicand(MPYF_mpd),.multiplier(MPYF_mpr),.signed_MPD(MPYF_MPD_sign),.signed_MPR(MPYF_MPR_sign));
MPY8x8 MPY_K(.csa_a(MPYK_csa_a),.csa_b(MPYK_csa_b),.multiplicand(MPYK_mpd),.multiplier(MPYK_mpr),.signed_MPD(MPYK_MPD_sign),.signed_MPR(MPYK_MPR_sign));



wire	[15:0] MPYG_cla_ina, MPYG_cla_inb;

assign MPYG_cla_ina = MPYG_csa_a;
assign MPYG_cla_inb = MPYG_csa_b;

wire	CLA16_G_g, CLA16_G_p, MPYG_ci;
assign MPYG_ci = 1'b0;

wire dangle_g_nodeJ, dangle_p_nodeJ; 
wire dangle_g_nodeF, dangle_p_nodeF; 
wire dangle_g_nodeK, dangle_p_nodeK; 



fcla16 CLA16_G(
.Sum(MPYG_o[15:0]),
.A(MPYG_cla_ina[15:0]),
.B(MPYG_cla_inb[15:0]), 
.G(CLA16_G_g),
.P(CLA16_G_p),
.Cin(MPYG_ci)
);



fcla16 CLA16_J(
.Sum(MPYJ_o[15:0]),
.A(MPYJ_csa_a[15:0]),
.B(MPYJ_csa_b[15:0]), 
.Cin(1'b0),
.G(dangle_g_nodeJ),
.P(dangle_p_nodeJ)
);



fcla16 CLA16_F(
.Sum(MPYF_o[15:0]),
.A(MPYF_csa_a[15:0]),
.B(MPYF_csa_b[15:0]), 
.Cin(1'b0),
.G(dangle_g_nodeF),
.P(dangle_p_nodeF)
);


fcla16 CLA16_K(
.Sum(MPYK_o[15:0]),
.A(MPYK_csa_a[15:0]),
.B(MPYK_csa_b[15:0]), 
.Cin(1'b0),
.G(dangle_g_nodeK), 
.P(dangle_p_nodeK)
);



always @(posedge clk or posedge IHRST)
begin
  if (IHRST)
    MPYF_oreg <= 0;		//#1 0;
  else
    MPYF_oreg <= MPYF_o; 	//#1 MPYF_o;
end

always @(posedge clk or posedge IHRST)
begin
  if (IHRST)
    MPYJ_oreg <=0; 		//#1 0;
  else if (MPY_8X8_MODE)
    MPYJ_oreg <=MPYJ_oreg;	//#1 MPYJ_oreg;
  else
    MPYJ_oreg <=MPYJ_o;  	//#1 MPYJ_o;
end

always @(posedge clk or posedge ILRST)
begin
  if (ILRST)
    MPYK_oreg <=0; 		//#1 0;
  else if (MPY_8X8_MODE)
    MPYK_oreg <=MPYK_oreg; 	//#1 MPYK_oreg;
  else
    MPYK_oreg <=MPYK_o; 	//#1 MPYK_o;
end

always @(posedge clk or posedge ILRST)
begin
  if (ILRST)
    MPYG_oreg <= 0; 		//#1 0;
  else
    MPYG_oreg <= MPYG_o; 	//#1 MPYG_o;
end

 assign MPYG_out = GSEL ? MPYG_oreg : MPYG_o;
 assign MPYJ_out = JKSEL ? MPYJ_oreg : MPYJ_o;

 assign MPYF_out = JKSEL ? MPYF_oreg : MPYF_o;
 assign MPYK_out = FSEL ? MPYK_oreg : MPYK_o;

wire [23:0] csa_oc;
wire [23:0] csa_os;
wire MPYJK_g_b;
assign MPYJK_g_b = ~MPYJK_g;

assign csa_os[23] = MPYJK_p ^ MPYF_out[15];
assign csa_oc[23] = ~(MPYJK_g_b & ~(MPYJK_p & MPYF_out[15]));
assign csa_os[22] = MPYJK_p ^ MPYF_out[14];
assign csa_oc[22] = ~(MPYJK_g_b & ~(MPYJK_p & MPYF_out[14]));
assign csa_os[21] = MPYJK_p ^ MPYF_out[13];
assign csa_oc[21] = ~(MPYJK_g_b & ~(MPYJK_p & MPYF_out[13]));
assign csa_os[20] = MPYJK_p ^ MPYF_out[12];
assign csa_oc[20] = ~(MPYJK_g_b & ~(MPYJK_p & MPYF_out[12]));
assign csa_os[19] = MPYJK_p ^ MPYF_out[11];
assign csa_oc[19] = ~(MPYJK_g_b & ~(MPYJK_p & MPYF_out[11]));
assign csa_os[18] = MPYJK_p ^ MPYF_out[10];
assign csa_oc[18] = ~(MPYJK_g_b & ~(MPYJK_p & MPYF_out[10]));
assign csa_os[17] = MPYJK_p ^ MPYF_out[9];
assign csa_oc[17] = ~(MPYJK_g_b & ~(MPYJK_p & MPYF_out[9]));
assign csa_os[16] = MPYJK_p ^ MPYF_out[8];
assign csa_oc[16] = ~(MPYJK_g_b & ~(MPYJK_p & MPYF_out[8]));

fa FA1_R00C15(.Cout(csa_oc[15]), .Sum(csa_os[15]), .A(MPYJ_out[15]), .B(MPYK_out[15]), .C(MPYF_out[7]));
fa FA1_R00C14(.Cout(csa_oc[14]), .Sum(csa_os[14]), .A(MPYJ_out[14]), .B(MPYK_out[14]), .C(MPYF_out[6]));
fa FA1_R00C13(.Cout(csa_oc[13]), .Sum(csa_os[13]), .A(MPYJ_out[13]), .B(MPYK_out[13]), .C(MPYF_out[5]));
fa FA1_R00C12(.Cout(csa_oc[12]), .Sum(csa_os[12]), .A(MPYJ_out[12]), .B(MPYK_out[12]), .C(MPYF_out[4]));
fa FA1_R00C11(.Cout(csa_oc[11]), .Sum(csa_os[11]), .A(MPYJ_out[11]), .B(MPYK_out[11]), .C(MPYF_out[3]));
fa FA1_R00C10(.Cout(csa_oc[10]), .Sum(csa_os[10]), .A(MPYJ_out[10]), .B(MPYK_out[10]), .C(MPYF_out[2]));
fa FA1_R00C09(.Cout(csa_oc[9]),  .Sum(csa_os[9]),  .A(MPYJ_out[9]),  .B(MPYK_out[9]),  .C(MPYF_out[1]));
fa FA1_R00C08(.Cout(csa_oc[8]),  .Sum(csa_os[8]),  .A(MPYJ_out[8]),  .B(MPYK_out[8]),  .C(MPYF_out[0]));

fa FA1_R00C07(.Cout(csa_oc[7]), .Sum(csa_os[7]), .A(MPYG_out[15]), .B(MPYJ_out[7]), .C(MPYK_out[7]));
fa FA1_R00C06(.Cout(csa_oc[6]), .Sum(csa_os[6]), .A(MPYG_out[14]), .B(MPYJ_out[6]), .C(MPYK_out[6]));
fa FA1_R00C05(.Cout(csa_oc[5]), .Sum(csa_os[5]), .A(MPYG_out[13]), .B(MPYJ_out[5]), .C(MPYK_out[5]));
fa FA1_R00C04(.Cout(csa_oc[4]), .Sum(csa_os[4]), .A(MPYG_out[12]), .B(MPYJ_out[4]), .C(MPYK_out[4]));
fa FA1_R00C03(.Cout(csa_oc[3]), .Sum(csa_os[3]), .A(MPYG_out[11]), .B(MPYJ_out[3]), .C(MPYK_out[3]));
fa FA1_R00C02(.Cout(csa_oc[2]), .Sum(csa_os[2]), .A(MPYG_out[10]), .B(MPYJ_out[2]), .C(MPYK_out[2]));
fa FA1_R00C01(.Cout(csa_oc[1]), .Sum(csa_os[1]), .A(MPYG_out[9]),  .B(MPYJ_out[1]), .C(MPYK_out[1]));
fa FA1_R00C00(.Cout(csa_oc[0]), .Sum(csa_os[0]), .A(MPYG_out[8]),  .B(MPYJ_out[0]), .C(MPYK_out[0]));


wire 	[23:0] cla_ina;
wire 	[23:0] cla_inb;

wire 	[23:0] cla_o;
wire	cla24_g0, cla24_p0;
wire	cla24_g1, cla24_p1;

wire	cla24_cin, cla24_16_cout;

assign cla_ina = csa_os;
assign cla_inb = {csa_oc[22:0],1'b0};
assign cla24_cin = 1'b0 ;


fcla16 CLA24_16(
.Sum(cla_o[15:0]),
.G(cla24_g0),
.P(cla24_p0), 
.A(cla_ina[15:0]),
.B(cla_inb[15:0]), 
.Cin(cla24_cin)
);
assign cla24_16_cout = ~(~cla24_g0 & ~(cla24_p0 & cla24_cin));



fcla8 CLA24_8(
.Sum(cla_o[23:16]),
.G(cla24_g1),
.P(cla24_p1), 
.A(cla_ina[23:16]),
.B(cla_inb[23:16]), 
.Cin(cla24_16_cout)
);

reg 	[31:0]mpy16_reg;

always @(posedge clk or posedge ILRST)
begin
  if (ILRST)
    mpy16_reg <= 0; 		//#1 0;
  else if (MPY_8X8_MODE)
    mpy16_reg <=  mpy16_reg; 	//#1 mpy16_reg;
  else
    mpy16_reg <={cla_o,MPYG_out[7:0]}; 	//#1 {cla_o,MPYG_out[7:0]};
end

assign O_16X16[31:0] = HSEL ? mpy16_reg : {cla_o,MPYG_out[7:0]};

assign OH_8X8 = MPYF_out[15:0];
assign OL_8X8 = MPYG_out[15:0];

endmodule // MPY16x16


//////////////////////////////////////////////////////////////////////////////////

`timescale 1ns / 1ps

module MULT_ACCUM(
    DIRECT_INPUT,
    MULT_INPUT,
    MULT_8x8,
    MULT_16x16,
	ADDSUB,
	CLK,
    CICAS,
    CI,
	SIGNEXTIN,
	SIGNEXTOUT,
    LDA,
    RST,
    ENA,
    COCAS,
    CO,
    O,
	OUTMUX_SEL,
	CARRYMUX_SEL,
	ADDER_A_IN_SEL,
	ADDER_B_IN_SEL
    );
	
    input [15:0] DIRECT_INPUT;
    input [15:0] MULT_INPUT;
    input [15:0] MULT_8x8;
    input [15:0] MULT_16x16;
    input ADDSUB;
    input CLK;
    input CICAS;
    input CI;
    input SIGNEXTIN;
    output SIGNEXTOUT;
    input LDA;
    input RST;
    input ENA;
    output COCAS;
    output CO;
    output [15:0] O;
	input [1:0] OUTMUX_SEL;
	input [1:0] CARRYMUX_SEL;
	input ADDER_A_IN_SEL;
	input [1:0] ADDER_B_IN_SEL;

	
	 wire [15:0] ADDER_LOAD_MUX ;
	 wire [15:0] ACCUMULATOR_REG ;
	 wire [15:0] ADDER_SUM ;
	 wire [15:0] ADDER_A_INPUT_MUX ;
	 wire [15:0] ADDER_B_INPUT_MUX ;
	 wire ADDER_CI ;
	 
	 assign SIGNEXTOUT = ADDER_B_INPUT_MUX[15];
	 

OUT_MUX_4 OUTPUT_MULTIPLEXER_TOP (
    .ADDER_COMBINATORIAL (ADDER_LOAD_MUX),
	 .ACCUM_REGISTER(ACCUMULATOR_REG) ,
	 .MULT_8x8(MULT_8x8) ,
	 .MULT_16x16(MULT_16x16),
	 .SELM(OUTMUX_SEL[1:0]) ,
	 .OUT(O)  
	 ) ;
	 
ACCUM_REG ACCUM_REG_TOP (
	.D(ADDER_LOAD_MUX) ,
	.Q(ACCUMULATOR_REG) ,
	.ENA(ENA) ,
	.CLK(CLK) ,
	.RST(RST)
	);
	
ACCUM_ADDER ACCUM_ADDER_TOP(
   .A(ADDER_A_INPUT_MUX) ,
   .B(ADDER_B_INPUT_MUX) ,
	.ADDSUB(ADDSUB) ,
	.CI(ADDER_CI) ,
	.SUM(ADDER_SUM) ,
	.COCAS(COCAS) ,
	.CO(CO)
	);	

LOAD_ADD_MUX LOAD_ADD_TOP (
   .ADDER(ADDER_SUM) ,
	.LOAD_DATA(DIRECT_INPUT) ,
	.LOAD(LDA),
	.OUT(ADDER_LOAD_MUX)
   );
	
ADDER_A_IN_MUX ADDER_A_IN_MUX_TOP (
   .ACCUMULATOR_REG(ACCUMULATOR_REG),
	.DIRECT_INPUT(DIRECT_INPUT) ,
	.SELM(ADDER_A_IN_SEL) ,
	.ADDER_A_MUX(ADDER_A_INPUT_MUX)
   );

ADDER_B_IN_MUX ADDER_B_IN_MUX_TOP (
   .MULT_INPUT(MULT_INPUT) ,
	.MULT_8x8(MULT_8x8) ,
	.MULT_16x16(MULT_16x16) ,
	.SIGNEXTIN(SIGNEXTIN) ,
	.SELM(ADDER_B_IN_SEL[1:0]) ,
	.ADDER_B_MUX(ADDER_B_INPUT_MUX)
	);	

CARRY_IN_MUX CARRY_IN_MUX_TOP (
	.CICAS(CICAS),
	.CI(CI),
	.CARRYMUX_SEL(CARRYMUX_SEL[1:0]),
	.ADDER_CI(ADDER_CI)
	);
	
endmodule

///////////////////////////////////////////////////////////////////////////////////
`timescale 1ns / 1ps

module OUT_MUX_4 (
    ADDER_COMBINATORIAL ,
	ACCUM_REGISTER ,
	MULT_8x8 ,
	MULT_16x16 ,
	SELM ,
	OUT  
	 ) ;

    input [15:0] ADDER_COMBINATORIAL ;
	input [15:0] ACCUM_REGISTER ;
	input [15:0] MULT_8x8 ;
	input [15:0] MULT_16x16 ;
	input [1:0] SELM ;
	output [15:0] OUT;  
	reg [15:0] OUT;  
	 
 
always @(SELM or ADDER_COMBINATORIAL or ACCUM_REGISTER or MULT_8x8 or MULT_16x16)
      case (SELM[1:0])
         2'b00: OUT = ADDER_COMBINATORIAL ; // Combinatorial output
         2'b01: OUT = ACCUM_REGISTER ; // Accumulator register output
         2'b10: OUT = MULT_8x8;  // MULT_8x8
         2'b11: OUT = MULT_16x16;  // MULT_16x16
      endcase	 

endmodule


///////////////////////////////////////////////////////////////////////

`timescale 1ns / 1ps

module ACCUM_REG (
	D ,
	Q ,
	ENA ,
	CLK ,
	RST
	);

	input [15:0] D ;
	output [15:0] Q;
	reg [15:0] Q;
	input ENA ;
	input CLK ;
	input RST;
	
	always @(posedge CLK or posedge RST)
      if (RST) // Syncronous reset overrides all other controls
				Q <= 16'h0 ;
		else
			if(ENA) // Update Q whenever LOAD or ENAble asserted
			    Q <=  D ; 	 //#1 D ;
			else
			    Q <= Q ;     //#1 Q ;
		
endmodule 


///////////////////////////////////////////////////////////////////////
`timescale 1ns / 1ps

module LOAD_ADD_MUX (
    ADDER ,
	LOAD_DATA ,
	LOAD,
	OUT
   );

	input [15:0] ADDER ;
	input [15:0] LOAD_DATA ;
	input LOAD;
	output [15:0] OUT;
   
	assign OUT = ( (LOAD) ? LOAD_DATA : ADDER ) ;
	
endmodule


///////////////////////////////////////////////////////////////////////
`timescale 1ns / 1ps

module ADDER_A_IN_MUX (
    ACCUMULATOR_REG ,
	DIRECT_INPUT ,
	SELM ,
	ADDER_A_MUX
   );
	
    input [15:0] ACCUMULATOR_REG ;
	input [15:0] DIRECT_INPUT ;
	input SELM ;
	output [15:0] ADDER_A_MUX;

	assign ADDER_A_MUX = ( (SELM) ? DIRECT_INPUT : ACCUMULATOR_REG ) ;

endmodule


///////////////////////////////////////////////////////////////////////
`timescale 1ns / 1ps

module ADDER_B_IN_MUX (
    MULT_INPUT ,
	MULT_8x8 ,
	MULT_16x16 ,
	SIGNEXTIN ,
	SELM ,
	ADDER_B_MUX
	);

    input [15:0] MULT_INPUT ;
	input [15:0] MULT_8x8 ;
	input [15:0] MULT_16x16 ;
	input SIGNEXTIN ;
	input [1:0] SELM ;
	output [15:0] ADDER_B_MUX;
	
//	wire [15:0] DIRECT_8x8_SELECT ;
//	assign DIRECT_8x8_SELECT = ( (SELM[0]) ? MULT_8x8   : MULT_INPUT) ;
//	assign ADDER_B_MUX       = ( (SELM[1:0]=2'b10) ? MULT_16x16 : DIRECT_8x8_SELECT) ;

	reg [15:0] ADDER_B_MUX;
	
always @(SELM or MULT_INPUT or MULT_8x8 or MULT_16x16 or SIGNEXTIN)
      case (SELM[1:0])
         2'b00: ADDER_B_MUX = MULT_INPUT ; 
         2'b01: ADDER_B_MUX = MULT_8x8 ; 
         2'b10: ADDER_B_MUX = MULT_16x16; 
         2'b11: ADDER_B_MUX = {16{SIGNEXTIN}}; 
      endcase	 
	
endmodule


///////////////////////////////////////////////////////////////////////

`timescale 1ns / 1ps
module CARRY_IN_MUX (
	CICAS,
	CI,
	CARRYMUX_SEL,
	ADDER_CI
	);
	
	input CICAS;
	input CI;
	input [1:0] CARRYMUX_SEL;
	output ADDER_CI;
	reg ADDER_CI;
	
always @(CARRYMUX_SEL or CICAS or CI)
      case (CARRYMUX_SEL[1:0])
         2'b00: ADDER_CI = 0 ; 
         2'b01: ADDER_CI = 1 ; 
         2'b10: ADDER_CI = CICAS; 
         2'b11: ADDER_CI = CI; 
      endcase	 

endmodule
	
//////////////////////////////////////////////////////////////////////////////////

`timescale 1ns / 1ps

module ACCUM_ADDER (
	A ,
	B ,
	ADDSUB ,
	CI ,
	SUM ,
	COCAS ,
	CO
	);
//parameter A_width =16;
input [15:0] A ;
input [15:0] B ;
input ADDSUB ;
input CI ;
output [15:0] SUM ;
output COCAS, CO;

wire	CLA16_g, CLA16_p;
reg		CO;

wire [15:0] CLA16_SUM;
reg	[15:0] CLA16_A, SUM;
integer j;

always@(ADDSUB or COCAS or A or CLA16_SUM)
begin
	if (ADDSUB)
		begin
		   CO = ~COCAS;
           for (j=0; j<=15; j=j+1)
			begin
			 CLA16_A[j] = ~A[j];
			 SUM[j] = ~CLA16_SUM[j];
			end 
		end   
		else
		begin
		   CO = COCAS;
		   CLA16_A[15:0] = A[15:0];
		   SUM[15:0] = CLA16_SUM[15:0];
		end
end

fcla16 CLA16_ADDER(
.Sum(CLA16_SUM[15:0]),
.A(CLA16_A[15:0]),
.B(B[15:0]), 
.G(CLA16_g),
.P(CLA16_p),
.Cin(CI)
);
assign COCAS= ~(~CLA16_g & ~(CLA16_p & CI));


endmodule


///////////////////////////////////////////////////////////////////////

`timescale 1ns / 1ps

module ha (Cout, Sum, A, B);
input A, B;
output Cout, Sum;

assign Cout = A & B;
assign Sum  = A ^ B;

endmodule // ha

///////////////////////////////////////////////////////////////////////

`timescale 1ns / 1ps
module fa (Cout, Sum, A, B, C);
input A, B, C;
output Cout, Sum;

//assign Cout = ((A&B) | (B&C) |(A&C));

assign Cout = ~(~(A&B) & ~(B&C) & ~(A&C));
assign Sum  = A^B^C;

endmodule // fa

///////////////////////////////////////////////////////////////////////

`timescale 1ns / 1ps

module mpfa (g_b, p,Sum, A, B, Cin);
input A, B, Cin;
output g_b, p, Sum;


assign g_b = ~(A & B);
assign p = A ^ B;

assign Sum  = p ^ Cin;

endmodule // mpfa

///////////////////////////////////////////////////////////////////////

`timescale 1ns / 1ps

module mclg4 (cout, g_o, p_o, g_b, p, cin);
input [3:0] g_b, p;
input cin;
output [3:0] cout;
output g_o, p_o;

wire	s1, s2, s3, s4, s5, s6,s7,s8,s9;

wire  [2:0] g;
assign g[0] =~g_b[0];
assign g[1] =~g_b[1];
assign g[2] =~g_b[2];

assign s1 = ~(p[0] & cin);
assign cout[1] =~(g_b[0] & s1);

assign s2 = ~(p[1] & g[0]);
assign s3 = ~(p[1] & p[0] & cin);
assign cout[2] =~(g_b[1] & s2 & s3);

assign s4 = ~(p[2] & g[1]);
assign s5 = ~(p[2] & p[1] & g[0]);
assign s6 = ~(p[2] & p[1] & p[0] & cin);
assign cout[3] =~(g_b[2] & s4 & s5 & s6);

assign s7 =~(p[3] & g[2]);
assign s8 =~(p[3] & p[2] & g[1]);
assign s9 =~(p[3] & p[2] & p[1] & g[0]);
assign g_o =~(g_b[3] & s7 & s8 & s9);

assign p_o =(p[3] & p[2] & p[1] & p[0]);

endmodule // mclg4

///////////////////////////////////////////////////////////////////////

`timescale 1ns / 1ps

module mclg16 (cout, g_o, p_o, g, p, cin);
input [3:0] g, p;
input cin;
output [3:0] cout;
output g_o, p_o;

wire	s1, s2, s3, s4, s5, s6, s7,s8,s9;

assign s1 = ~(p[0] & cin);
assign cout[1] =~(~g[0] & s1);

assign s2 = ~(p[1] & g[0]);
assign s3 = ~(p[1] & p[0] & cin);
assign cout[2] =~(~g[1] & s2 & s3);

assign s4 = ~(p[2] & g[1]);
assign s5 = ~(p[2] & p[1] & g[0]);
assign s6 = ~(p[2] & p[1] & p[0] & cin);
assign cout[3] =~(~g[2] & s4 & s5 & s6);

assign s7 =~(p[3] & g[2]);
assign s8 =~(p[3] & p[2] & g[1]);
assign s9 =~(p[3] & p[2] & p[1] & g[0]);
assign g_o =~(~g[3] & s7 & s8 & s9);

assign p_o =(p[3] & p[2] & p[1] & p[0]);

endmodule // mclg16
///////////////////////////////////////////////////////////////////////


`timescale 1ns / 1ps
module fcla16 (Sum, G, P, A, B, Cin);
input [15:0] A, B;
input Cin;
output [15:0] Sum;
output G, P;
wire	[15:0] gtemp1_b;
wire	[15:0] ptemp1;
wire	[15:0] ctemp1;
wire	[3:0] ctemp2;

wire	[3:0] gouta, pouta;
mpfa r01 (.g_b(gtemp1_b[0]), .p(ptemp1[0]), .Sum(Sum[0]), .A(A[0]), .B(B[0]), .Cin(Cin));
mpfa r02 (.g_b(gtemp1_b[1]), .p(ptemp1[1]), .Sum(Sum[1]), .A(A[1]), .B(B[1]), .Cin(ctemp1[1]));
mpfa r03 (.g_b(gtemp1_b[2]), .p(ptemp1[2]), .Sum(Sum[2]), .A(A[2]), .B(B[2]), .Cin(ctemp1[2]));
mpfa r04 (.g_b(gtemp1_b[3]), .p(ptemp1[3]), .Sum(Sum[3]), .A(A[3]), .B(B[3]), .Cin(ctemp1[3]));
mclg4 b1 (.cout(ctemp1[3:0]), .g_o(gouta[0]), .p_o(pouta[0]), .g_b(gtemp1_b[3:0]), .p(ptemp1[3:0]), .cin(Cin));

mpfa r05 (.g_b(gtemp1_b[4]), .p(ptemp1[4]), .Sum(Sum[4]), .A(A[4]), .B(B[4]), .Cin(ctemp2[1]));
mpfa r06 (.g_b(gtemp1_b[5]), .p(ptemp1[5]), .Sum(Sum[5]), .A(A[5]), .B(B[5]), .Cin(ctemp1[5]));
mpfa r07 (.g_b(gtemp1_b[6]), .p(ptemp1[6]), .Sum(Sum[6]), .A(A[6]), .B(B[6]), .Cin(ctemp1[6]));
mpfa r08 (.g_b(gtemp1_b[7]), .p(ptemp1[7]), .Sum(Sum[7]), .A(A[7]), .B(B[7]), .Cin(ctemp1[7]));
mclg4 b2 (.cout(ctemp1[7:4]), .g_o(gouta[1]), .p_o(pouta[1]), .g_b(gtemp1_b[7:4]), .p(ptemp1[7:4]), .cin(ctemp2[1]));

mpfa r09 (.g_b(gtemp1_b[8]), .p(ptemp1[8]), .Sum(Sum[8]), .A(A[8]), .B(B[8]), .Cin(ctemp2[2]));
mpfa r10 (.g_b(gtemp1_b[9]), .p(ptemp1[9]), .Sum(Sum[9]), .A(A[9]), .B(B[9]), .Cin(ctemp1[9]));
mpfa r11 (.g_b(gtemp1_b[10]), .p(ptemp1[10]), .Sum(Sum[10]), .A(A[10]), .B(B[10]), .Cin(ctemp1[10]));
mpfa r12 (.g_b(gtemp1_b[11]), .p(ptemp1[11]), .Sum(Sum[11]), .A(A[11]), .B(B[11]), .Cin(ctemp1[11]));
mclg4 b3 (.cout(ctemp1[11:8]), .g_o(gouta[2]), .p_o(pouta[2]), .g_b(gtemp1_b[11:8]), .p(ptemp1[11:8]), .cin(ctemp2[2]));

mpfa r13 (.g_b(gtemp1_b[12]), .p(ptemp1[12]), .Sum(Sum[12]), .A(A[12]), .B(B[12]), .Cin(ctemp2[3]));
mpfa r14 (.g_b(gtemp1_b[13]), .p(ptemp1[13]), .Sum(Sum[13]), .A(A[13]), .B(B[13]), .Cin(ctemp1[13]));
mpfa r15 (.g_b(gtemp1_b[14]), .p(ptemp1[14]), .Sum(Sum[14]), .A(A[14]), .B(B[14]), .Cin(ctemp1[14]));
mpfa r16 (.g_b(gtemp1_b[15]), .p(ptemp1[15]), .Sum(Sum[15]), .A(A[15]), .B(B[15]), .Cin(ctemp1[15]));
mclg4 b4 (.cout(ctemp1[15:12]), .g_o(gouta[3]), .p_o(pouta[3]), .g_b(gtemp1_b[15:12]), .p(ptemp1[15:12]), .cin(ctemp2[3]));

mclg16 b5 (.cout(ctemp2), .g_o(G), .p_o(P), .g(gouta), .p(pouta), .cin(Cin));
endmodule // fcla16


///////////////////////////////////////////////////////////////////////

`timescale 1ns / 1ps

module fcla8 (Sum, G, P, A, B, Cin);
input [7:0] A, B;
input Cin;
output [7:0] Sum;
output G, P;
wire	[7:0] gtemp1;
wire	[7:0] ptemp1;
wire	[7:0] ctemp1;
wire	 ctemp2;

wire	[1:0] gouta, pouta;

mpfa r01 (.g_b(gtemp1[0]), .p(ptemp1[0]), .Sum(Sum[0]), .A(A[0]), .B(B[0]), .Cin(Cin));
mpfa r02 (.g_b(gtemp1[1]), .p(ptemp1[1]), .Sum(Sum[1]), .A(A[1]), .B(B[1]), .Cin(ctemp1[1]));
mpfa r03 (.g_b(gtemp1[2]), .p(ptemp1[2]), .Sum(Sum[2]), .A(A[2]), .B(B[2]), .Cin(ctemp1[2]));
mpfa r04 (.g_b(gtemp1[3]), .p(ptemp1[3]), .Sum(Sum[3]), .A(A[3]), .B(B[3]), .Cin(ctemp1[3]));
mclg4 b1 (.cout(ctemp1[3:0]), .g_o(gouta[0]), .p_o(pouta[0]), .g_b(gtemp1[3:0]), .p(ptemp1[3:0]), .cin(Cin));

mpfa r05 (.g_b(gtemp1[4]), .p(ptemp1[4]), .Sum(Sum[4]), .A(A[4]), .B(B[4]), .Cin(ctemp2));
mpfa r06 (.g_b(gtemp1[5]), .p(ptemp1[5]), .Sum(Sum[5]), .A(A[5]), .B(B[5]), .Cin(ctemp1[5]));
mpfa r07 (.g_b(gtemp1[6]), .p(ptemp1[6]), .Sum(Sum[6]), .A(A[6]), .B(B[6]), .Cin(ctemp1[6]));
mpfa r08 (.g_b(gtemp1[7]), .p(ptemp1[7]), .Sum(Sum[7]), .A(A[7]), .B(B[7]), .Cin(ctemp1[7]));
mclg4 b2 (.cout(ctemp1[7:4]), .g_o(gouta[1]), .p_o(pouta[1]), .g_b(gtemp1[7:4]), .p(ptemp1[7:4]), .cin(ctemp2));

assign ctemp2=~(~gouta[0] & ~(pouta[0] & Cin));

assign G = ~(~gouta[1] & ~(pouta[1] & gouta[0]));
assign P = pouta[1] & pouta[0];

endmodule // fcla8


//////////////////////////////////////////////////////////////////////////////// 

`timescale 1ns / 1ps

module REG_BYPASS_MUX(D, Q, ENA, CLK, RST, SELM);

parameter DATA_WIDTH = 16 ;

input  [DATA_WIDTH - 1 : 0] D ;
output [DATA_WIDTH - 1 : 0] Q ;
input  ENA ;
input  CLK ;
input  RST ;
input  SELM ;

reg    [DATA_WIDTH - 1 : 0] REG_INTERNAL ;

assign Q = ( (SELM) ? REG_INTERNAL : D ) ;

always @ (posedge CLK or posedge RST)
begin
	if (RST)
		REG_INTERNAL <= #1 0 ;
	else if (ENA)
	    REG_INTERNAL <= #1 D ;
	else 
	    REG_INTERNAL <= #1 REG_INTERNAL ;
end

endmodule



//----------------------------------------------//
//---  SB_IO_DLY Synthesis Primitive -----------// 
//---------------------------------------------// 

`timescale 10ps/1ps

module SB_IO_DLY (
	PACKAGE_PIN, 
	LATCH_INPUT_VALUE, 
	CLOCK_ENABLE, 
	INPUT_CLK, 
	OUTPUT_CLK, 
	OUTPUT_ENABLE, 
	D_OUT_1, 
	D_OUT_0, 
	D_IN_1, 
	D_IN_0,
	SCLK,
	SDI,
	C_R_SEL,
	SDO
 );


parameter NEG_TRIGGER 	= 1'b0; 	   // When set to 1'b1 the polarity of all FFs in the IO is set work at falling edge, default is rising edge Flops
parameter PIN_TYPE      = 6'b000000;       // The required package pin type must be set when io_macro is instantiated.
parameter PULLUP 	= 1'b0;	
parameter IO_STANDARD 	= "SB_LVCMOS";     
parameter INDELAY_VAL   = 6'b000000;       // Set input  line delay value 
parameter OUTDELAY_VAL  = 6'b000000;       // Set output line delay value 


inout 	PACKAGE_PIN; 		//' User's package pin - 'PAD' output
input 	CLOCK_ENABLE;    	// Clock enables in & out clocks
input 	LATCH_INPUT_VALUE;    	// Input Latch data control
input	INPUT_CLK;   		// Input clock
input 	OUTPUT_CLK;  		// Output clock


output 	D_IN_1;    		// Data to Core from PAD     - input 1   (ddrin1)
output	D_IN_0;    		// Data to Core from PAD     - input 0   (ddrin0)

input 	D_OUT_1;  		// Data to PAD from core - output 1 (ddrout1)
input 	D_OUT_0;  		// Data to PAD from core - output 0 (ddrout0)  
input 	OUTPUT_ENABLE;   	// Ouput-Enable 

input  SCLK;			// Delay serial register clock  
input  SDI;                     // Serial data input to serial delay registers  
input  C_R_SEL;                 //'0' selects IN/OUT static delay parameters, '1' selects serial register data 
output SDO;                     // Serial data out from serial registers 


//------------- Main Body of verilog ----------------------------------------------------
wire inclk_, outclk_;
wire inclk, outclk;
reg INCLKE_sync, OUTCLKE_sync;

assign (weak0, weak1) CLOCK_ENABLE =1'b1 ;
assign inclk_ = (INPUT_CLK ^ NEG_TRIGGER); // change the input clock phase
assign outclk_ = (OUTPUT_CLK ^ NEG_TRIGGER); // change the output clock phase
//assign inclk = (inclk_ & CLOCK_ENABLE);
//assign outclk = (outclk_ & CLOCK_ENABLE);

//////// CLKEN sync ///////
always@(inclk_ or CLOCK_ENABLE)
begin 
    if(~inclk_)
	INCLKE_sync = CLOCK_ENABLE; 
end

always@(outclk_ or CLOCK_ENABLE)
begin 
   if(~outclk_) 	
	OUTCLKE_sync = CLOCK_ENABLE; 
end

assign inclk = (inclk_ & INCLKE_sync);
assign outclk = (outclk_ & OUTCLKE_sync);

wire bs_en;   //Boundary scan enable
wire shift;   //Boundary scan shift
wire tclk;    //Boundary scan clock
wire update;  //Boundary scan update
wire sdi;     //Boundary scan serial data in
wire mode;    //Boundary scan mode
wire hiz_b;   //Boundary scan tristate control
wire sdo;     //Boundary scan serial data out

//wire rstio; disabled as this a power on only signal   	//Normal Input reset
assign  bs_en = 1'b0;	//Boundary scan enable
assign  shift = 1'b0;	//Boundary scan shift
assign  tclk = 1'b0;	//Boundary scan clock
assign  update = 1'b0;	//Boundary scan update
assign  sdi = 1'b0;	//Boundary scan serial data in
assign  mode = 1'b0;	//Boundary scan mode
assign  hiz_b = 1'b1;	//Boundary scan Tristate control
  
wire padoen, padout, padin;
wire padinout_delayed; 
assign PACKAGE_PIN = (~padoen) ? padinout_delayed : 1'bz;
assign padin = PACKAGE_PIN ;

wire hold, oepin;							  
assign hold = LATCH_INPUT_VALUE;
assign oepin = OUTPUT_ENABLE;
 
 preio_physical preiophysical_i (	//original names unchanged
 	.hold(hold),
	.rstio(1'b0),			//Disabled as this is power on only.
	.bs_en(bs_en),
	.shift(shift),
	.tclk(tclk),
	.inclk(inclk),
	.outclk(outclk),
	.update(update),
	.oepin(oepin),
	.sdi(sdi),
	.mode(mode),
	.hiz_b(hiz_b),
	.sdo(sdo),
	.dout1(D_IN_1),
	.dout0(D_IN_0),
	.ddr1(D_OUT_1),
	.ddr0(D_OUT_0),
	.padin(padinout_delayed),
	.padout(padout),
	.padoen(padoen),
	.cbit(PIN_TYPE)
	);

   inoutdly64 iodly64_i ( 
	// dynamic delay test logic thru sdi , sdo pins disabled // 
	.sclk(),
        .serialreg_rst(),
        .sdi(),
        .c_r_sel(),
        .in_datain(padin),
        .out_datain(padout),
        .delay_direction(padoen),
        .delayed_dataout(padinout_delayed),
        .sdo()
	); 
   defparam iodly64_i.INDELAY  =INDELAY_VAL; 
   defparam iodly64_i.OUTDELAY =OUTDELAY_VAL; 
    	        

`ifdef TIMINGCHECK
specify
   // tp,tCQ to din0/din1 
   (PACKAGE_PIN *> D_IN_0) = (1.0, 1.0);
   (INPUT_CLK *> D_IN_0) = (1.0, 1.0);
   (INPUT_CLK *> D_IN_1) = (1.0, 1.0);
   (LATCH_INPUT_VALUE *> D_IN_0) = (1.0, 1.0);
   //tp,tCQ to PP  
   (D_OUT_0 *> PACKAGE_PIN) = (1.0, 1.0);
   (OUTPUT_ENABLE *> PACKAGE_PIN) = (1.0, 1.0);
   (OUTPUT_CLK *> PACKAGE_PIN) = (1.0, 1.0);
   //CE-INCLK 	
   $setup(posedge CLOCK_ENABLE, posedge INPUT_CLK, 1.0);
   $setup(negedge CLOCK_ENABLE, posedge INPUT_CLK, 1.0);
   $hold(posedge INPUT_CLK, posedge CLOCK_ENABLE, 1.0);
   $hold(posedge INPUT_CLK, negedge CLOCK_ENABLE, 1.0);
   //CE-OUTCLK
   $setup(posedge CLOCK_ENABLE, posedge OUTPUT_CLK, 1.0);
   $setup(negedge CLOCK_ENABLE, posedge OUTPUT_CLK, 1.0);
   $hold(posedge OUTPUT_CLK, posedge CLOCK_ENABLE, 1.0);
   $hold(posedge OUTPUT_CLK, negedge CLOCK_ENABLE, 1.0);
   //setup/hold wrt posedge iclk (DIN0 reg)  
   $setup(posedge PACKAGE_PIN, posedge INPUT_CLK, 1.0);
   $setup(negedge PACKAGE_PIN, posedge INPUT_CLK, 1.0);
   $hold(posedge INPUT_CLK, posedge PACKAGE_PIN, 1.0);
   $hold(posedge INPUT_CLK, negedge PACKAGE_PIN, 1.0);
   //setup/hold wrt negedge iclk (DIN1 reg)  
   $setup(posedge PACKAGE_PIN, negedge INPUT_CLK, 1.0);
   $setup(negedge PACKAGE_PIN, negedge INPUT_CLK, 1.0);
   $hold(negedge INPUT_CLK, posedge PACKAGE_PIN, 1.0);
   $hold(negedge INPUT_CLK, negedge PACKAGE_PIN, 1.0);
   // setup/hold wrt to posedge oclk (DOUT0 reg) 
   $setup(posedge D_OUT_0, posedge OUTPUT_CLK, 1.0);
   $setup(negedge D_OUT_0, posedge OUTPUT_CLK, 1.0);
   $hold(posedge OUTPUT_CLK, posedge D_OUT_0, 1.0);
   $hold(posedge OUTPUT_CLK, negedge D_OUT_0, 1.0);
   // setup/hold wrt to negedge oclk (DOUT1 reg) 
   $setup(posedge D_OUT_1, negedge OUTPUT_CLK, 1.0);
   $setup(negedge D_OUT_1, negedge OUTPUT_CLK, 1.0);
   $hold(negedge OUTPUT_CLK, posedge D_OUT_1, 1.0);
   $hold(negedge OUTPUT_CLK, negedge D_OUT_1, 1.0);
   // setup/hold wrt to posedge oclk (OE reg)
   $setup(posedge OUTPUT_ENABLE, posedge OUTPUT_CLK, 1.0);
   $setup(negedge OUTPUT_ENABLE, posedge OUTPUT_CLK, 1.0);
   $hold(posedge OUTPUT_CLK, posedge OUTPUT_ENABLE, 1.0);
   $hold(posedge OUTPUT_CLK, negedge OUTPUT_ENABLE, 1.0);
endspecify
`endif

endmodule


//----------------------------------------------------// 
//-----    64 TAP DELAY LOGIC ------------------------//
//----------------------------------------------------//

`timescale 1ps/1ps 	

module inoutdly64 (
		sclk,
		serialreg_rst,
		sdi,
		c_r_sel,
		in_datain, 
		out_datain, 
		delay_direction, 
		delayed_dataout,
		sdo 
);

parameter 	INDELAY  = 6'b000000;
parameter 	OUTDELAY = 6'b000000;

localparam	BUF_DELAY=100;	  	// 100ps +-25 ps 
localparam     	CBITS_DELAY ={OUTDELAY,INDELAY};  

input	sclk;		// shiftreg serial clock 
input	serialreg_rst; 	// delay register reset 
input	sdi;          	// serial data in 
input	c_r_sel; 	// Select Cbits or ShiftRegister Value for Delay    
input 	in_datain;  	// padin  data to delay tap 
input 	out_datain;      // padout data to delay tap 
input 	delay_direction;      // delay tap direction. 0 -Apply delay on output data to PAD, 1 -Apply delay on input data from PAD. 
			// delay_direction is controlled by oen of PRE_IO model.  
output	sdo;            // serial data out.
output	delayed_dataout;	// delayed data output   

reg  [11:0] cbits; 
reg  [11:0] serial_data;  
wire [5:0]  delay_sel; 
wire 	    data_in; 

wire [63:1] buf_y; 
reg         delayed_data; 

integer i; 

initial 
begin
 for(i=0 ; i<12 ; i=i+1) 
 begin 
  cbits[i]	=CBITS_DELAY[i]; 	// initialize cbits value 	
 end
 serial_data =12'b0; 
end 

// serial dynamic delay data  
always@(posedge sclk or posedge serialreg_rst) 
begin 
	if(serialreg_rst ==1'b1) 
		serial_data <= 12'b0; 
//	else  						// left shift 
//		serial_data <= {serial_data[10:0],sdi};
	else						// right shift 
		serial_data <= {sdi,serial_data[11:1]}; 
end
assign	sdo = serial_data[0]; 

// SDI, SDO dynamic delay test sections is not required. Delays are static and based on the in out delay parameters.  
//assign delay_sel = (delay_direction == 1'b0)?(c_r_sel ==1'b0)? cbits[11:6]:serial_data[11:6] : (c_r_sel ==1'b0)? cbits[5:0]:serial_data[5:0]; 

assign delay_sel = (delay_direction == 1'b0) ? OUTDELAY    : INDELAY; 
assign data_in   = (delay_direction == 1'b0) ? out_datain  : in_datain ; 

// 63 buf tap  
buf #BUF_DELAY  bufinst1 (buf_y[1],data_in );   
buf #BUF_DELAY  bufinst2 (buf_y[2],buf_y[1]);   
buf #BUF_DELAY  bufinst3 (buf_y[3],buf_y[2]);   
buf #BUF_DELAY  bufinst4 (buf_y[4],buf_y[3]);   
buf #BUF_DELAY  bufinst5 (buf_y[5],buf_y[4]);   
buf #BUF_DELAY  bufinst6 (buf_y[6],buf_y[5]);   
buf #BUF_DELAY  bufinst7 (buf_y[7],buf_y[6]);   
buf #BUF_DELAY  bufinst8 (buf_y[8],buf_y[7]);   
buf #BUF_DELAY  bufinst9 (buf_y[9],buf_y[8]);   
buf #BUF_DELAY  bufinst10 (buf_y[10],buf_y[9]); 

buf #BUF_DELAY  bufinst11 (buf_y[11],buf_y[10]);
buf #BUF_DELAY  bufinst12 (buf_y[12],buf_y[11]);
buf #BUF_DELAY  bufinst13 (buf_y[13],buf_y[12]);
buf #BUF_DELAY  bufinst14 (buf_y[14],buf_y[13]);
buf #BUF_DELAY  bufinst15 (buf_y[15],buf_y[14]);
buf #BUF_DELAY  bufinst16 (buf_y[16],buf_y[15]);
buf #BUF_DELAY  bufinst17 (buf_y[17],buf_y[16]); 
buf #BUF_DELAY  bufinst18 (buf_y[18],buf_y[17]); 
buf #BUF_DELAY  bufinst19 (buf_y[19],buf_y[18]); 
buf #BUF_DELAY  bufinst20 (buf_y[20],buf_y[19]); 

buf #BUF_DELAY  bufinst21 (buf_y[21],buf_y[20] );
buf #BUF_DELAY  bufinst22 (buf_y[22],buf_y[21]); 
buf #BUF_DELAY  bufinst23 (buf_y[23],buf_y[22]); 
buf #BUF_DELAY  bufinst24 (buf_y[24],buf_y[23]); 
buf #BUF_DELAY  bufinst25 (buf_y[25],buf_y[24]); 
buf #BUF_DELAY  bufinst26 (buf_y[26],buf_y[25]); 
buf #BUF_DELAY  bufinst27 (buf_y[27],buf_y[26]); 
buf #BUF_DELAY  bufinst28 (buf_y[28],buf_y[27]); 
buf #BUF_DELAY  bufinst29 (buf_y[29],buf_y[28]); 
buf #BUF_DELAY  bufinst30 (buf_y[30],buf_y[29]); 

buf #BUF_DELAY  bufinst31 (buf_y[31],buf_y[30]); 
buf #BUF_DELAY  bufinst32 (buf_y[32],buf_y[31]); 
buf #BUF_DELAY  bufinst33 (buf_y[33],buf_y[32]); 
buf #BUF_DELAY  bufinst34 (buf_y[34],buf_y[33]); 
buf #BUF_DELAY  bufinst35 (buf_y[35],buf_y[34]); 
buf #BUF_DELAY  bufinst36 (buf_y[36],buf_y[35]); 
buf #BUF_DELAY  bufinst37 (buf_y[37],buf_y[36]); 
buf #BUF_DELAY  bufinst38 (buf_y[38],buf_y[37]); 
buf #BUF_DELAY  bufinst39 (buf_y[39],buf_y[38]); 
buf #BUF_DELAY  bufinst40 (buf_y[40],buf_y[39]); 

buf #BUF_DELAY  bufinst41 (buf_y[41],buf_y[40]); 
buf #BUF_DELAY  bufinst42 (buf_y[42],buf_y[41]); 
buf #BUF_DELAY  bufinst43 (buf_y[43],buf_y[42]); 
buf #BUF_DELAY  bufinst44 (buf_y[44],buf_y[43]); 
buf #BUF_DELAY  bufinst45 (buf_y[45],buf_y[44]); 
buf #BUF_DELAY  bufinst46 (buf_y[46],buf_y[45]); 
buf #BUF_DELAY  bufinst47 (buf_y[47],buf_y[46]); 
buf #BUF_DELAY  bufinst48 (buf_y[48],buf_y[47]); 
buf #BUF_DELAY  bufinst49 (buf_y[49],buf_y[48]); 
buf #BUF_DELAY  bufinst50 (buf_y[50],buf_y[49]); 

buf #BUF_DELAY  bufinst51 (buf_y[51],buf_y[50]); 
buf #BUF_DELAY  bufinst52 (buf_y[52],buf_y[51]); 
buf #BUF_DELAY  bufinst53 (buf_y[53],buf_y[52]); 
buf #BUF_DELAY  bufinst54 (buf_y[54],buf_y[53]); 
buf #BUF_DELAY  bufinst55 (buf_y[55],buf_y[54]); 
buf #BUF_DELAY  bufinst56 (buf_y[56],buf_y[55]); 
buf #BUF_DELAY  bufinst57 (buf_y[57],buf_y[56]); 
buf #BUF_DELAY  bufinst58 (buf_y[58],buf_y[57]); 
buf #BUF_DELAY  bufinst59 (buf_y[59],buf_y[58]); 
buf #BUF_DELAY  bufinst60 (buf_y[60],buf_y[59]); 

buf #BUF_DELAY  bufinst61 (buf_y[61],buf_y[60]); 
buf #BUF_DELAY  bufinst62 (buf_y[62],buf_y[61]);   
buf #BUF_DELAY  bufinst63 (buf_y[63],buf_y[62]);   

// delay_sel mux 
always @*
begin 
	case(delay_sel) 
	6'd0: delayed_data  = data_in;   
	6'd1: delayed_data  = buf_y[1];    
	6'd2: delayed_data  = buf_y[2];  
	6'd3: delayed_data  = buf_y[3];
	6'd4: delayed_data  = buf_y[4];
	6'd5: delayed_data  = buf_y[5];
	6'd6: delayed_data  = buf_y[6];
	6'd7: delayed_data  = buf_y[7];
	6'd8: delayed_data  = buf_y[8];
	6'd9: delayed_data  = buf_y[9];
	6'd10: delayed_data = buf_y[10 ];

	6'd11: delayed_data = buf_y[11];
	6'd12: delayed_data = buf_y[12];
	6'd13: delayed_data = buf_y[13];
	6'd14: delayed_data = buf_y[14];
	6'd15: delayed_data = buf_y[15];
	6'd16: delayed_data = buf_y[16];
	6'd17: delayed_data = buf_y[17];
	6'd18: delayed_data = buf_y[18];
	6'd19: delayed_data = buf_y[19];
	6'd20: delayed_data = buf_y[20];

	6'd21: delayed_data = buf_y[21];
	6'd22: delayed_data = buf_y[22];
	6'd23: delayed_data = buf_y[23];
	6'd24: delayed_data = buf_y[24];
	6'd25: delayed_data = buf_y[25];
	6'd26: delayed_data = buf_y[26];
	6'd27: delayed_data = buf_y[27];
	6'd28: delayed_data = buf_y[28];
	6'd29: delayed_data = buf_y[29];
	6'd30: delayed_data = buf_y[30];

	6'd31: delayed_data = buf_y[31];
	6'd32: delayed_data = buf_y[32];
	6'd33: delayed_data = buf_y[33];
	6'd34: delayed_data = buf_y[34];
	6'd35: delayed_data = buf_y[35];
	6'd36: delayed_data = buf_y[36];
	6'd37: delayed_data = buf_y[37];
	6'd38: delayed_data = buf_y[38];
	6'd39: delayed_data = buf_y[39];
	6'd40: delayed_data = buf_y[40];

	6'd41: delayed_data = buf_y[41];
	6'd42: delayed_data = buf_y[42];
	6'd43: delayed_data = buf_y[43];
	6'd44: delayed_data = buf_y[44];
	6'd45: delayed_data = buf_y[45];
	6'd46: delayed_data = buf_y[46];
	6'd47: delayed_data = buf_y[47];
	6'd48: delayed_data = buf_y[48];
	6'd49: delayed_data = buf_y[49];
	6'd50: delayed_data = buf_y[50];

	6'd51: delayed_data = buf_y[51];
	6'd52: delayed_data = buf_y[52];
	6'd53: delayed_data = buf_y[53];
	6'd54: delayed_data = buf_y[54];
	6'd55: delayed_data = buf_y[55];
	6'd56: delayed_data = buf_y[56];
	6'd57: delayed_data = buf_y[57];
	6'd58: delayed_data = buf_y[58];
	6'd59: delayed_data = buf_y[59];
	6'd60: delayed_data = buf_y[60];

	6'd61: delayed_data = buf_y[61];
	6'd62: delayed_data = buf_y[62];
	6'd63: delayed_data = buf_y[63];
	endcase
end 

assign delayed_dataout = delayed_data ; 

endmodule

//---------------------------------------------------// 
//---- SB_MIPI_TX_4LANE Synthesis Primitive ---------//
//---------------------------------------------------//
`timescale 1ps/1ps
module    SB_MIPI_TX_4LANE (
//Common Interface Pins
input 		PU,
input		LBEN,
input 	[1:0]	ROUTCAL,
input 		ENPDESER,
input       	PDCKG,

// DATA0 Interface pins
inout		DP0,
inout		DN0,
input 		D0OPMODE,
input 		D0DTXLPP,
input 		D0DTXLPN,
input  		D0TXLPEN,
output 		D0DRXLPP,
output  	D0DRXLPN,
input 		D0RXLPEN,
output 		D0DCDP,
output		D0DCDN,
input 		D0CDEN,
input  		D0TXHSPD,
input 		D0TXHSEN,
input    [7:0]  D0HSTXDATA,
input  		D0HSSEREN,
input 		D0RXHSEN,
input  		D0HSDESEREN,
output 	 [7:0]	D0HSRXDATA,
output 		D0HSBYTECLKD,
output 		D0SYNC,
output 		D0ERRSYNC,
output      	D0HSBYTECLKSNOSYNC,
// DATA1 Interface pins
inout		DP1,
inout		DN1,
input 		D1DTXLPP,
input 		D1DTXLPN,
input  		D1TXLPEN,
output 		D1DRXLPP,
output  	D1DRXLPN,
input 		D1RXLPEN,
output 		D1DCDP,
output		D1DCDN,
input 		D1CDEN,
input  		D1TXHSPD,
input 		D1TXHSEN, 
input    [7:0]  D1HSTXDATA,
input  		D1HSSEREN,
input 		D1RXHSEN,
input  		D1HSDESEREN,
output 	 [7:0]	D1HSRXDATA,
output 		D1SYNC,
output 		D1ERRSYNC,
output 		D1NOSYNC,
// DATA2 Interface pins
inout		DP2,
inout		DN2,
input 		D2DTXLPP,
input 		D2DTXLPN,
input  		D2TXLPEN,
output 		D2DRXLPP,
output  	D2DRXLPN,
input 		D2RXLPEN,
output 		D2DCDP,
output		D2DCDN,
input 		D2CDEN,
input  		D2TXHSPD,
input 		D2TXHSEN, 
input    [7:0] 	D2HSTXDATA,
input  		D2HSSEREN,
input 		D2RXHSEN,
input  		D2HSDESEREN,
output 	 [7:0]	D2HSRXDATA,
output 		D2SYNC,
output 		D2ERRSYNC,
output 		D2NOSYNC,
// DATA3 Interface pins
inout		DP3,
inout		DN3,
input 		D3DTXLPP,
input 		D3DTXLPN,
input  		D3TXLPEN,
output 		D3DRXLPP,
output  	D3DRXLPN,
input 		D3RXLPEN,
output 		D3DCDP,
output		D3DCDN,
input 		D3CDEN,
input  		D3TXHSPD,
input 		D3TXHSEN, 
input    [7:0] 	D3HSTXDATA,
input  		D3HSSEREN,
input 		D3RXHSEN,
input  		D3HSDESEREN,
output 	 [7:0]	D3HSRXDATA,
output 		D3SYNC,
output 		D3ERRSYNC,
output 		D3NOSYNC,
// CLOCK Interface pins
inout		CKP,
inout		CKN,
input 		CLKDTXLPP,
input 		CLKDTXLPN,
input  		CLKTXLPEN,
output  	CLKDRXLPP,
output  	CLKDRXLPN,
input  		CLKRXLPEN,
input  		CLKTXHSPD,
input 		CLKTXHSEN,
input       	CLKTXHSGATE,
input  		CLKRXHSEN,
output      	CLKHSBYTE,
// Universal MIPI PLL Interface pins
input 		PLLPU,
input 		PLLREF,
output 		PLLLOCK,
//Universal MIPI PLL Serial Configuration Register Interface pins
input 		PLLCFGSRDI,
input 		PLLCFGSRRESET,
input 		PLLCFGSRCLK,
output 		PLLCFGSRDO
);
//parameter PLLCFG_DEFAULT = 20'h00000;
parameter DIVR = 5'b11111;   //Ref Clk divider
parameter DIVF = 8'b11110000; // Feedback divider
parameter DIVQ = 2'b00;       // VCO divider
parameter TEST_MODE = 1'b0;
parameter TEST_BITS = 4'b1001;

wire BITCLK_int; 

X1082T001 u_mipi_txrx_analog(
	// Power and Grd Pins 
	.VDDA(1'b1),
	.VSSA(1'b0),
	.VDD(1'b1),
	.VSS(1'b0),
	.DVSS(1'b0),
	//Common Interface Pins
	.BITCLK(BITCLK_int) ,
	.PD(~PU),
	.LB_EN(LBEN),
	.ROUT_CAL(ROUTCAL),
	.ENP_DESER(ENPDESER),
	.PDCKG(PDCKG),
	// DATA0 Interface pins
	.DP0(DP0),
	.DN0(DN0),
	.D0_OPMODE(D0OPMODE), 		// Input from digital to indicate mode of operation TX or RX
	.D0_DTXLPP(D0DTXLPP),
	.D0_DTXLPN(D0DTXLPN),
	.D0_TXLPEN(D0TXLPEN),
	.D0_DRXLPP(D0DRXLPP),
	.D0_DRXLPN(D0DRXLPN),
	.D0_RXLPEN(D0RXLPEN),
	.D0_DCDP(D0DCDP),
	.D0_DCDN(D0DCDN),
	.D0_CDEN(D0CDEN),
	.D0_TXHSPD(D0TXHSPD),
	.D0_TXHSEN(D0TXHSEN),
	.D0_HSTX_DATA(D0HSTXDATA),
	.D0_HS_SER_EN(D0HSSEREN),
	.D0_RXHSEN(D0RXHSEN),
	.D0_HS_DESER_EN(D0HSDESEREN),
	.D0_HSRX_DATA(D0HSRXDATA),
	.D0_HS_BYTE_CLKD(D0HSBYTECLKD), // Byteclk output from Lane0 deserializer
	.D0_SYNC(D0SYNC),
	.D0_ERRSYNC(D0ERRSYNC),
	.D0_HS_BYTE_CLKS_NOSYNC(D0HSBYTECLKSNOSYNC), // This output will be D0_NOSYNC or D0_HS_BYTE_CLKS based on D0_OPMODE
	// DATA1 Interface pins
	.DP1(DP1),
	.DN1(DN1),
	.D1_DTXLPP(D1DTXLPP),
	.D1_DTXLPN(D1DTXLPN),
	.D1_TXLPEN(D1TXLPEN),
	.D1_DRXLPP(D1DRXLPP),
	.D1_DRXLPN(D1DRXLPN),
	.D1_RXLPEN(D1RXLPEN),
	.D1_DCDP(D1DCDP),
	.D1_DCDN(D1DCDN),
	.D1_CDEN(D1CDEN),
	.D1_TXHSPD(D1TXHSPD),
	.D1_TXHSEN(D1TXHSEN),
	.D1_HSTX_DATA(D1HSTXDATA),
	.D1_HS_SER_EN(D1HSSEREN),
	.D1_RXHSEN(D1RXHSEN),
	.D1_HS_DESER_EN(D1HSDESEREN),
	.D1_HSRX_DATA(D1HSRXDATA),
	.D1_SYNC(D1SYNC),
	.D1_ERRSYNC(D1ERRSYNC),
	.D1_NOSYNC(D1NOSYNC),
	// DATA2 Interface pins
	.DP2(DP2),
	.DN2(DN2),
	.D2_DTXLPP(D2DTXLPP),
	.D2_DTXLPN(D2DTXLPN),
	.D2_TXLPEN(D2TXLPEN),
	.D2_DRXLPP(D2DRXLPP),
	.D2_DRXLPN(D2DRXLPN),
	.D2_RXLPEN(D2RXLPEN),
	.D2_DCDP(D2DCDP),
	.D2_DCDN(D2DCDN),
	.D2_CDEN(D2CDEN),
	.D2_TXHSPD(D2TXHSPD),
	.D2_TXHSEN(D2TXHSEN),
	.D2_HSTX_DATA(D2HSTXDATA),
	.D2_HS_SER_EN(D2HSSEREN),
	.D2_RXHSEN(D2RXHSEN),
	.D2_HS_DESER_EN(D2HSDESEREN),
	.D2_HSRX_DATA(D2HSRXDATA),
	.D2_SYNC(D2SYNC),
	.D2_ERRSYNC(D2ERRSYNC),
	.D2_NOSYNC(D2NOSYNC),
	// DATA3 Interface pins
	.DP3(DP3),
	.DN3(DN3),
	.D3_DTXLPP(D3DTXLPP),
	.D3_DTXLPN(D3DTXLPN),
	.D3_TXLPEN(D3TXLPEN),
	.D3_DRXLPP(D3DRXLPP),
	.D3_DRXLPN(D3DRXLPN),
	.D3_RXLPEN(D3RXLPEN),
	.D3_DCDP(D3DCDP),
	.D3_DCDN(D3DCDN),
	.D3_CDEN(D3CDEN),
	.D3_TXHSPD(D3TXHSPD),
	.D3_TXHSEN(D3TXHSEN),
	.D3_HSTX_DATA(D3HSTXDATA),
	.D3_HS_SER_EN(D3HSSEREN),
	.D3_RXHSEN(D3RXHSEN),
	.D3_HS_DESER_EN(D3HSDESEREN),
	.D3_HSRX_DATA(D3HSRXDATA),
	.D3_SYNC(D3SYNC),
	.D3_ERRSYNC(D3ERRSYNC),
	.D3_NOSYNC(D3NOSYNC),
	// CLOCK Interface pins
	.CKP(CKP),
	.CKN(CKN),
	.CLK_DTXLPP(CLKDTXLPP),
	.CLK_DTXLPN(CLKDTXLPN),
	.CLK_TXLPEN(CLKTXLPEN),
	.CLK_DRXLPP(CLKDRXLPP),
	.CLK_DRXLPN(CLKDRXLPN),
	.CLK_RXLPEN(CLKRXLPEN),
	.CLK_TXHSPD(CLKTXHSPD),
	.CLK_TXHSEN(CLKTXHSEN),
	.CLK_TXHSGATE(CLKTXHSGATE),
	.CLK_RXHSEN(CLKRXHSEN),
	.CLK_HS_BYTE(CLKHSBYTE)
);

X109T001 u_mipi_txpll_analog (
	.VDDA(1'b1),
	.VSSA(1'b0),
	.VDD(1'b1),
	.VSS(1'b0),
	.PD(~PLLPU), 
	.TST(4'b0),       
	.CN(DIVR),
	.CM(DIVF),
	.CO(DIVQ),
	.CLKREF(PLLREF),
	.OUTP(BITCLK_int),
	.OUTN(),
	.LOCK(PLLLOCK)	
 );


`ifdef TIMINGCHECK
specify
   // --- TX conf timing paths  ------// 	
   // Data0 lane tp & tCQ (TX conf) 	
   (D0DTXLPP *> DP0) = (1.0, 1.0); 
   (D0DTXLPN *> DN0) = (1.0, 1.0);
   (DP1      *> DP0) = (1.0, 1.0);  //tx-rx loop back  
   (DP1      *> DN0) = (1.0, 1.0);  //tx-rx loop back  
   (PLLREF   *> DP0) = (1.0, 1.0);   
   (PLLREF   *> DN0) = (1.0, 1.0); 
   (PLLREF   *> D0HSBYTECLKSNOSYNC) = (1.0,1.0); 	 
   // Data1 lane tp & tCQ (TX conf) 	
   (D1DTXLPP *> DP1) = (1.0, 1.0); 
   (D1DTXLPN *> DN1) = (1.0, 1.0);
   (DP0      *> DP1) = (1.0, 1.0);  //tx-rx loop back   
   (DP0      *> DN1) = (1.0, 1.0);  //tx-rx loop back   
   (PLLREF   *> DP1) = (1.0, 1.0);   
   (PLLREF   *> DN1) = (1.0, 1.0); 
   // Data2 lane tp & tCQ (TX conf) 	
   (D2DTXLPP *> DP2) = (1.0, 1.0); 
   (D2DTXLPN *> DN2) = (1.0, 1.0);
   (DP3      *> DP2) = (1.0, 1.0);  //tx-rx loop back   
   (DP3      *> DN2) = (1.0, 1.0);  //tx-rx loop back   
   (PLLREF   *> DP2) = (1.0, 1.0);   
   (PLLREF   *> DN2) = (1.0, 1.0); 
   // Data3 lane tp & tCQ (TX conf) 	
   (D3DTXLPP *> DP3) = (1.0, 1.0); 
   (D3DTXLPN *> DN3) = (1.0, 1.0);
   (DP2      *> DP3) = (1.0, 1.0);  //tx-rx loop back   
   (DP2      *> DN3) = (1.0, 1.0);  //tx-rx loop back   
   (PLLREF   *> DP3) = (1.0, 1.0);   
   (PLLREF   *> DN3) = (1.0, 1.0);   	
   //Clk Lane tp & tCQ (TX conf) 			 
   (CLKDTXLPP *> CKP) = (1.0,1.0);
   (CLKDTXLPN *> CKN) = (1.0,1.0);
   (PLLREF    *> CKP) = (1.0,1.0);
   (PLLREF    *> CKN) = (1.0,1.0);  
   // Data0 Lane setup-hold checks (TX conf)
   $setup(posedge D0HSTXDATA[0], posedge PLLREF, 1.0);
   $setup(negedge D0HSTXDATA[0], posedge PLLREF, 1.0);
   $hold (posedge PLLREF, posedge D0HSTXDATA[0], 1.0);
   $hold (posedge PLLREF, negedge D0HSTXDATA[0], 1.0);   
   $setup(posedge D0HSTXDATA[1], posedge PLLREF, 1.0);
   $setup(negedge D0HSTXDATA[1], posedge PLLREF, 1.0);
   $hold (posedge PLLREF, posedge D0HSTXDATA[1], 1.0);
   $hold (posedge PLLREF, negedge D0HSTXDATA[1], 1.0);   
   $setup(posedge D0HSTXDATA[2], posedge PLLREF, 1.0);
   $setup(negedge D0HSTXDATA[2], posedge PLLREF, 1.0);
   $hold (posedge PLLREF, posedge D0HSTXDATA[2], 1.0);
   $hold (posedge PLLREF, negedge D0HSTXDATA[2], 1.0);   
   $setup(posedge D0HSTXDATA[3], posedge PLLREF, 1.0);
   $setup(negedge D0HSTXDATA[3], posedge PLLREF, 1.0);
   $hold (posedge PLLREF, posedge D0HSTXDATA[3], 1.0);
   $hold (posedge PLLREF, negedge D0HSTXDATA[3], 1.0);   
   $setup(posedge D0HSTXDATA[4], posedge PLLREF, 1.0);
   $setup(negedge D0HSTXDATA[4], posedge PLLREF, 1.0);
   $hold (posedge PLLREF, posedge D0HSTXDATA[4], 1.0);
   $hold (posedge PLLREF, negedge D0HSTXDATA[4], 1.0);   
   $setup(posedge D0HSTXDATA[5], posedge PLLREF, 1.0);
   $setup(negedge D0HSTXDATA[5], posedge PLLREF, 1.0);
   $hold (posedge PLLREF, posedge D0HSTXDATA[5], 1.0);
   $hold (posedge PLLREF, negedge D0HSTXDATA[5], 1.0);   
   $setup(posedge D0HSTXDATA[6], posedge PLLREF, 1.0);
   $setup(negedge D0HSTXDATA[6], posedge PLLREF, 1.0);
   $hold (posedge PLLREF, posedge D0HSTXDATA[6], 1.0);
   $hold (posedge PLLREF, negedge D0HSTXDATA[6], 1.0);   
   $setup(posedge D0HSTXDATA[7], posedge PLLREF, 1.0);
   $setup(negedge D0HSTXDATA[7], posedge PLLREF, 1.0);
   $hold (posedge PLLREF, posedge D0HSTXDATA[7], 1.0);
   $hold (posedge PLLREF, negedge D0HSTXDATA[7], 1.0);   
   // Data1 Lane setup-hold checks (TX conf)
   $setup(posedge D1HSTXDATA[0], posedge PLLREF, 1.0);
   $setup(negedge D1HSTXDATA[0], posedge PLLREF, 1.0);
   $hold (posedge PLLREF, posedge D1HSTXDATA[0], 1.0);
   $hold (posedge PLLREF, negedge D1HSTXDATA[0], 1.0);   
   $setup(posedge D1HSTXDATA[1], posedge PLLREF, 1.0);
   $setup(negedge D1HSTXDATA[1], posedge PLLREF, 1.0);
   $hold (posedge PLLREF, posedge D1HSTXDATA[1], 1.0);
   $hold (posedge PLLREF, negedge D1HSTXDATA[1], 1.0);   
   $setup(posedge D1HSTXDATA[2], posedge PLLREF, 1.0);
   $setup(negedge D1HSTXDATA[2], posedge PLLREF, 1.0);
   $hold (posedge PLLREF, posedge D1HSTXDATA[2], 1.0);
   $hold (posedge PLLREF, negedge D1HSTXDATA[2], 1.0);   
   $setup(posedge D1HSTXDATA[3], posedge PLLREF, 1.0);
   $setup(negedge D1HSTXDATA[3], posedge PLLREF, 1.0);
   $hold (posedge PLLREF, posedge D1HSTXDATA[3], 1.0);
   $hold (posedge PLLREF, negedge D1HSTXDATA[3], 1.0);   
   $setup(posedge D1HSTXDATA[4], posedge PLLREF, 1.0);
   $setup(negedge D1HSTXDATA[4], posedge PLLREF, 1.0);
   $hold (posedge PLLREF, posedge D1HSTXDATA[4], 1.0);
   $hold (posedge PLLREF, negedge D1HSTXDATA[4], 1.0);   
   $setup(posedge D1HSTXDATA[5], posedge PLLREF, 1.0);
   $setup(negedge D1HSTXDATA[5], posedge PLLREF, 1.0);
   $hold (posedge PLLREF, posedge D1HSTXDATA[5], 1.0);
   $hold (posedge PLLREF, negedge D1HSTXDATA[5], 1.0);   
   $setup(posedge D1HSTXDATA[6], posedge PLLREF, 1.0);
   $setup(negedge D1HSTXDATA[6], posedge PLLREF, 1.0);
   $hold (posedge PLLREF, posedge D1HSTXDATA[6], 1.0);
   $hold (posedge PLLREF, negedge D1HSTXDATA[6], 1.0);   
   $setup(posedge D1HSTXDATA[7], posedge PLLREF, 1.0);
   $setup(negedge D1HSTXDATA[7], posedge PLLREF, 1.0);
   $hold (posedge PLLREF, posedge D1HSTXDATA[7], 1.0);
   $hold (posedge PLLREF, negedge D1HSTXDATA[7], 1.0);   
   // Data2 Lane setup-hold checks (TX conf)
   $setup(posedge D2HSTXDATA[0], posedge PLLREF, 1.0);
   $setup(negedge D2HSTXDATA[0], posedge PLLREF, 1.0);
   $hold (posedge PLLREF, posedge D2HSTXDATA[0], 1.0);
   $hold (posedge PLLREF, negedge D2HSTXDATA[0], 1.0);   
   $setup(posedge D2HSTXDATA[1], posedge PLLREF, 1.0);
   $setup(negedge D2HSTXDATA[1], posedge PLLREF, 1.0);
   $hold (posedge PLLREF, posedge D2HSTXDATA[1], 1.0);
   $hold (posedge PLLREF, negedge D2HSTXDATA[1], 1.0);   
   $setup(posedge D2HSTXDATA[2], posedge PLLREF, 1.0);
   $setup(negedge D2HSTXDATA[2], posedge PLLREF, 1.0);
   $hold (posedge PLLREF, posedge D2HSTXDATA[2], 1.0);
   $hold (posedge PLLREF, negedge D2HSTXDATA[2], 1.0);   
   $setup(posedge D2HSTXDATA[3], posedge PLLREF, 1.0);
   $setup(negedge D2HSTXDATA[3], posedge PLLREF, 1.0);
   $hold (posedge PLLREF, posedge D2HSTXDATA[3], 1.0);
   $hold (posedge PLLREF, negedge D2HSTXDATA[3], 1.0);   
   $setup(posedge D2HSTXDATA[4], posedge PLLREF, 1.0);
   $setup(negedge D2HSTXDATA[4], posedge PLLREF, 1.0);
   $hold (posedge PLLREF, posedge D2HSTXDATA[4], 1.0);
   $hold (posedge PLLREF, negedge D2HSTXDATA[4], 1.0);   
   $setup(posedge D2HSTXDATA[5], posedge PLLREF, 1.0);
   $setup(negedge D2HSTXDATA[5], posedge PLLREF, 1.0);
   $hold (posedge PLLREF, posedge D2HSTXDATA[5], 1.0);
   $hold (posedge PLLREF, negedge D2HSTXDATA[5], 1.0);   
   $setup(posedge D2HSTXDATA[6], posedge PLLREF, 1.0);
   $setup(negedge D2HSTXDATA[6], posedge PLLREF, 1.0);
   $hold (posedge PLLREF, posedge D2HSTXDATA[6], 1.0);
   $hold (posedge PLLREF, negedge D2HSTXDATA[6], 1.0);   
   $setup(posedge D2HSTXDATA[7], posedge PLLREF, 1.0);
   $setup(negedge D2HSTXDATA[7], posedge PLLREF, 1.0);
   $hold (posedge PLLREF, posedge D2HSTXDATA[7], 1.0);
   $hold (posedge PLLREF, negedge D2HSTXDATA[7], 1.0);   
   // Data3 Lane setup-hold checks (TX conf)
   $setup(posedge D3HSTXDATA[0], posedge PLLREF, 1.0);
   $setup(negedge D3HSTXDATA[0], posedge PLLREF, 1.0);
   $hold (posedge PLLREF, posedge D3HSTXDATA[0], 1.0);
   $hold (posedge PLLREF, negedge D3HSTXDATA[0], 1.0);   
   $setup(posedge D3HSTXDATA[1], posedge PLLREF, 1.0);
   $setup(negedge D3HSTXDATA[1], posedge PLLREF, 1.0);
   $hold (posedge PLLREF, posedge D3HSTXDATA[1], 1.0);
   $hold (posedge PLLREF, negedge D3HSTXDATA[1], 1.0);   
   $setup(posedge D3HSTXDATA[2], posedge PLLREF, 1.0);
   $setup(negedge D3HSTXDATA[2], posedge PLLREF, 1.0);
   $hold (posedge PLLREF, posedge D3HSTXDATA[2], 1.0);
   $hold (posedge PLLREF, negedge D3HSTXDATA[2], 1.0);   
   $setup(posedge D3HSTXDATA[3], posedge PLLREF, 1.0);
   $setup(negedge D3HSTXDATA[3], posedge PLLREF, 1.0);
   $hold (posedge PLLREF, posedge D3HSTXDATA[3], 1.0);
   $hold (posedge PLLREF, negedge D3HSTXDATA[3], 1.0);   
   $setup(posedge D3HSTXDATA[4], posedge PLLREF, 1.0);
   $setup(negedge D3HSTXDATA[4], posedge PLLREF, 1.0);
   $hold (posedge PLLREF, posedge D3HSTXDATA[4], 1.0);
   $hold (posedge PLLREF, negedge D3HSTXDATA[4], 1.0);   
   $setup(posedge D3HSTXDATA[5], posedge PLLREF, 1.0);
   $setup(negedge D3HSTXDATA[5], posedge PLLREF, 1.0);
   $hold (posedge PLLREF, posedge D3HSTXDATA[5], 1.0);
   $hold (posedge PLLREF, negedge D3HSTXDATA[5], 1.0);   
   $setup(posedge D3HSTXDATA[6], posedge PLLREF, 1.0);
   $setup(negedge D3HSTXDATA[6], posedge PLLREF, 1.0);
   $hold (posedge PLLREF, posedge D3HSTXDATA[6], 1.0);
   $hold (posedge PLLREF, negedge D3HSTXDATA[6], 1.0);   
   $setup(posedge D3HSTXDATA[7], posedge PLLREF, 1.0);
   $setup(negedge D3HSTXDATA[7], posedge PLLREF, 1.0);
   $hold (posedge PLLREF, posedge D3HSTXDATA[7], 1.0);
   $hold (posedge PLLREF, negedge D3HSTXDATA[7], 1.0);   

    // --- RX conf timing paths -------// 
    //Data0 Lane tp & tCQ (RX conf) 
   (DP0 *> D0DRXLPP) = (1.0, 1.0);
   (DN0 *> D0DRXLPN) = (1.0, 1.0);	
   (DP0 *> D0DCDP  ) = (1.0, 1.0);	  
   (DN0 *> D0DCDN  ) = (1.0, 1.0); 
   (CKP *> D0HSRXDATA[0]) = (1.0, 1.0);	
   (CKP *> D0HSRXDATA[1]) = (1.0, 1.0);	
   (CKP *> D0HSRXDATA[2]) = (1.0, 1.0);	
   (CKP *> D0HSRXDATA[3]) = (1.0, 1.0);	
   (CKP *> D0HSRXDATA[4]) = (1.0, 1.0);	
   (CKP *> D0HSRXDATA[5]) = (1.0, 1.0);	
   (CKP *> D0HSRXDATA[6]) = (1.0, 1.0);	
   (CKP *> D0HSRXDATA[7]) = (1.0, 1.0);	
   (CKP *> D0HSBYTECLKD ) = (1.0, 1.0);	 
    //Data1 Lane tp & tCQ  (RX conf)
   (DP1 *> D1DRXLPP) = (1.0, 1.0);
   (DN1 *> D1DRXLPN) = (1.0, 1.0);	
   (DP1 *> D1DCDP  ) = (1.0, 1.0);	  
   (DN1 *> D1DCDN  ) = (1.0, 1.0); 
   (CKP *> D1HSRXDATA[0]) = (1.0, 1.0);	
   (CKP *> D1HSRXDATA[1]) = (1.0, 1.0);	
   (CKP *> D1HSRXDATA[2]) = (1.0, 1.0);	
   (CKP *> D1HSRXDATA[3]) = (1.0, 1.0);	
   (CKP *> D1HSRXDATA[4]) = (1.0, 1.0);	
   (CKP *> D1HSRXDATA[5]) = (1.0, 1.0);	
   (CKP *> D1HSRXDATA[6]) = (1.0, 1.0);	
   (CKP *> D1HSRXDATA[7]) = (1.0, 1.0);	
    //Data2 Lane tp & tCQ (RX conf) 
   (DP2 *> D2DRXLPP) = (1.0, 1.0);
   (DN2 *> D2DRXLPN) = (1.0, 1.0);
   (DP2 *> D2DCDP  ) = (1.0, 1.0);	  
   (DN2 *> D2DCDN  ) = (1.0, 1.0); 
   (CKP *> D2HSRXDATA[0]) = (1.0, 1.0);	
   (CKP *> D2HSRXDATA[1]) = (1.0, 1.0);	
   (CKP *> D2HSRXDATA[2]) = (1.0, 1.0);	
   (CKP *> D2HSRXDATA[3]) = (1.0, 1.0);	
   (CKP *> D2HSRXDATA[4]) = (1.0, 1.0);	
   (CKP *> D2HSRXDATA[5]) = (1.0, 1.0);	
   (CKP *> D2HSRXDATA[6]) = (1.0, 1.0);	
   (CKP *> D2HSRXDATA[7]) = (1.0, 1.0);	
    //Data3 Lane tp & tCQ (RX conf) 
   (DP3 *> D3DRXLPP) = (1.0, 1.0);
   (DN3 *> D3DRXLPN) = (1.0, 1.0);	
   (DP3 *> D3DCDP  ) = (1.0, 1.0);	  
   (DN3 *> D3DCDN  ) = (1.0, 1.0); 
   (CKP *> D3HSRXDATA[0]) = (1.0, 1.0);	
   (CKP *> D3HSRXDATA[1]) = (1.0, 1.0);	
   (CKP *> D3HSRXDATA[2]) = (1.0, 1.0);	
   (CKP *> D3HSRXDATA[3]) = (1.0, 1.0);	
   (CKP *> D3HSRXDATA[4]) = (1.0, 1.0);	
   (CKP *> D3HSRXDATA[5]) = (1.0, 1.0);	
   (CKP *> D3HSRXDATA[6]) = (1.0, 1.0);	
   (CKP *> D3HSRXDATA[7]) = (1.0, 1.0);	
   //Clk Lane tp & tCQ (RX conf) 			  
   (CKP  *> CLKDRXLPP ) = (1.0, 1.0);
   (CKN  *> CLKDRXLPN ) = (1.0, 1.0);
   (CKP  *> CLKHSBYTE) = (1.0, 1.0);
   // Data0 Lane setup-hold checks (RX conf)
   $setup(posedge DP0, posedge CKP, 1.0);
   $setup(negedge DP0, posedge CKP, 1.0);
   $hold (posedge CKP, posedge DP0, 1.0);
   $hold (posedge CKP, negedge DP0, 1.0);   
   $setup(posedge DP0, negedge CKP, 1.0);
   $setup(negedge DP0, negedge CKP, 1.0);
   $hold (negedge CKP, posedge DP0, 1.0);
   $hold (negedge CKP, negedge DP0, 1.0);
   
   $setup(posedge DN0, posedge CKP, 1.0);
   $setup(negedge DN0, posedge CKP, 1.0);
   $hold (posedge CKP, posedge DN0, 1.0);
   $hold (posedge CKP, negedge DN0, 1.0);   
   $setup(posedge DN0, negedge CKP, 1.0);
   $setup(negedge DN0, negedge CKP, 1.0);
   $hold (negedge CKP, posedge DN0, 1.0);
   $hold (negedge CKP, negedge DN0, 1.0);
   // Data1 Lane setup-hold checks (RX conf) 
   $setup(posedge DP1, posedge CKP, 1.0);
   $setup(negedge DP1, posedge CKP, 1.0);
   $hold (posedge CKP, posedge DP1, 1.0);
   $hold (posedge CKP, negedge DP1, 1.0);   
   $setup(posedge DP1, negedge CKP, 1.0);
   $setup(negedge DP1, negedge CKP, 1.0);
   $hold (negedge CKP, posedge DP1, 1.0);
   $hold (negedge CKP, negedge DP1, 1.0);  
   
   $setup(posedge DN1, posedge CKP, 1.0);
   $setup(negedge DN1, posedge CKP, 1.0);
   $hold (posedge CKP, posedge DN1, 1.0);
   $hold (posedge CKP, negedge DN1, 1.0);   
   $setup(posedge DN1, negedge CKP, 1.0);
   $setup(negedge DN1, negedge CKP, 1.0);
   $hold (negedge CKP, posedge DN1, 1.0);
   $hold (negedge CKP, negedge DN1, 1.0);      
   // Data2 Lane setup-hold cheks (RX conf) 
   $setup(posedge DP2, posedge CKP, 1.0);
   $setup(negedge DP2, posedge CKP, 1.0);
   $hold (posedge CKP, posedge DP2, 1.0);
   $hold (posedge CKP, negedge DP2, 1.0);   
   $setup(posedge DP2, negedge CKP, 1.0);
   $setup(negedge DP2, negedge CKP, 1.0);
   $hold (negedge CKP, posedge DP2, 1.0);
   $hold (negedge CKP, negedge DP2, 1.0);
   
   $setup(posedge DN2, posedge CKP, 1.0);
   $setup(negedge DN2, posedge CKP, 1.0);
   $hold (posedge CKP, posedge DN2, 1.0);
   $hold (posedge CKP, negedge DN2, 1.0);   
   $setup(posedge DN2, negedge CKP, 1.0);
   $setup(negedge DN2, negedge CKP, 1.0);
   $hold (negedge CKP, posedge DN2, 1.0);
   $hold (negedge CKP, negedge DN2, 1.0);
   // Data3 Lane setup-hold cheks (RX conf)
   $setup(posedge DP3, posedge CKP, 1.0);
   $setup(negedge DP3, posedge CKP, 1.0);
   $hold (posedge CKP, posedge DP3, 1.0);
   $hold (posedge CKP, negedge DP3, 1.0);   
   $setup(posedge DP3, negedge CKP, 1.0);
   $setup(negedge DP3, negedge CKP, 1.0);
   $hold (negedge CKP, posedge DP3, 1.0);
   $hold (negedge CKP, negedge DP3, 1.0);
   
   $setup(posedge DN3, posedge CKP, 1.0);
   $setup(negedge DN3, posedge CKP, 1.0);
   $hold (posedge CKP, posedge DN3, 1.0);
   $hold (posedge CKP, negedge DN3, 1.0);   
   $setup(posedge DN3, negedge CKP, 1.0);
   $setup(negedge DN3, negedge CKP, 1.0);
   $hold (negedge CKP, posedge DN3, 1.0);
   $hold (negedge CKP, negedge DN3, 1.0);
endspecify
`endif   



endmodule //SB_MIPI_TX_4LANE



//-----------------------------------------------------------------------------------------------------//
//              	---  ICE40MH - 16K Block RAM Primitives  -----  
// Front End Primitives :  
//	# SB_RAM1024x16		# SB_RAM1024x16NR  	# SB_RAM1024x16NW	# SB_RAM1024x16NRNW
//	# SB_RAM2048x8		# SB_RAM2048x8NR	# SB_RAM2048x8NW	# SB_RAM2048x8NRNW
//	# SB_RAM4096x4		# SB_RAM4096x4NR	# SB_RAM4096x4NW	# SB_RAM4096x4NRNW
//	# SB_RAM8192x2		# SB_RAM8192x2NR	# SB_RAM8192x2NW	# SB_RAM8192x2NRNW
// Back End Primitives  : 
//	# SB_RAM40_16K	   # SB_RAM40_16KNR 	# SB_RAM40_16KNW 	# SB_RAM40_16KNRNW
//-------------------------------------------------------------------------------------------------------//

//---------------------------------
//	-- SB_RAM1024x16 --
//---------------------------------
`timescale 1ps/1ps
module  SB_RAM1024x16 ( RDATA, RCLK, RCLKE, RE, RADDR, WCLK, WCLKE, WE, WADDR, MASK, WDATA );

output	[15:0]	RDATA;  
input         	RCLK;   
input           RCLKE; 
input           RE; 
input	[9:0]   RADDR; 
input           WCLK; 
input           WCLKE; 
input           WE; 
input 	[9:0]   WADDR; 
input	[15:0]	MASK; 
input 	[15:0]	WDATA; 

parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

// local Parameters
localparam			CLOCK_PERIOD = 200;	//
localparam 			DELAY	= (CLOCK_PERIOD/10);		// Clock-to-output delay. Zero
							// time delays can be confusing
							// and sometimes cause problems.
localparam 			BUS_WIDTH = 16;		// Width of RAM (number of bits)

localparam 			ADDRESS_BUS_SIZE = 10;	// Number of bits required to
							// represent the RAM address

localparam   ADDRESSABLE_SPACE  = 2**ADDRESS_BUS_SIZE;	// Decimal address range [2^Size:0]


// SIGNAL DECLARATIONS
wire			   	WCLK_g, RCLK_g;
reg 				WCLKE_sync, RCLKE_sync; 
assign (weak0, weak1) RCLKE =1'b1 ;
assign (weak0, weak1) RE =1'b0 ;
assign (weak0, weak1) WCLKE =1'b1 ;
assign (weak0, weak1) WE =1'b0 ;
reg	Memory	[BUS_WIDTH*ADDRESSABLE_SPACE-1:0];
// 
event Read_e, Write_e;

//////////////////// Collision detect begins here ///////////////////////////////
localparam 	TRUE = 1'b1;
localparam	FALSE = 1'b0;
reg 		Time_Collision_Detected = 1'b0;
wire		Address_Collision_Detected;

event Collision_e;

time COLLISION_TIME_WINDOW = (CLOCK_PERIOD/8); // This is an arbitray value, but is better than using an absolute 
						    // value, because the actual time window depends on the actual silicon 
						    // implementation. Thus the test is indicative of an Error and not
						    // guaranteed to be an error. Even so this is usefull.
time time_WCLK_RCLK, time_WCLK, time_RCLK;


//function reg Check_Timed_Window_Violation;
function	Check_Timed_Window_Violation;	
input T1, T2, Minimum_Time_Window;
time T1, T2;
time Minimum_Time_Window;
time Difference;	
	begin
		Difference = (T1 - T2);
		if (Difference < 0) Difference = -Difference;
		Check_Timed_Window_Violation = (Difference < Minimum_Time_Window);
	end
endfunction


initial begin
       time_WCLK = CLOCK_PERIOD;	// Arbitrary initialisation value, ensure no window collison error on first clock edge.
       time_RCLK = (CLOCK_PERIOD*8);	// Arbitrary initialisation difference value, ensure no collision error on first clock edge.					
end

integer	i,j;


initial	//	initialize ram_16k (1024 x 16) by init parameters, section by section
begin
	for	(i=0; i<=(256/BUS_WIDTH)-1; i=i+1)       
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)    
		begin 

			Memory[BUS_WIDTH*i+j]		=	INIT_0[BUS_WIDTH*i+j];
			Memory[256*1+BUS_WIDTH*i+j]	=	INIT_1[BUS_WIDTH*i+j];
			Memory[256*2+BUS_WIDTH*i+j]	=	INIT_2[BUS_WIDTH*i+j];
			Memory[256*3+BUS_WIDTH*i+j]	=	INIT_3[BUS_WIDTH*i+j];
			Memory[256*4+BUS_WIDTH*i+j]	=	INIT_4[BUS_WIDTH*i+j];
			Memory[256*5+BUS_WIDTH*i+j]	=	INIT_5[BUS_WIDTH*i+j];
			Memory[256*6+BUS_WIDTH*i+j]	=	INIT_6[BUS_WIDTH*i+j];
			Memory[256*7+BUS_WIDTH*i+j]	=	INIT_7[BUS_WIDTH*i+j];
			Memory[256*8+BUS_WIDTH*i+j]	=	INIT_8[BUS_WIDTH*i+j];
			Memory[256*9+BUS_WIDTH*i+j]	=	INIT_9[BUS_WIDTH*i+j];
			Memory[256*10+BUS_WIDTH*i+j]	=	INIT_A[BUS_WIDTH*i+j];
			Memory[256*11+BUS_WIDTH*i+j]	=	INIT_B[BUS_WIDTH*i+j];
			Memory[256*12+BUS_WIDTH*i+j]	=	INIT_C[BUS_WIDTH*i+j];
			Memory[256*13+BUS_WIDTH*i+j]	=	INIT_D[BUS_WIDTH*i+j];
			Memory[256*14+BUS_WIDTH*i+j]	=	INIT_E[BUS_WIDTH*i+j];
			Memory[256*15+BUS_WIDTH*i+j]	=	INIT_F[BUS_WIDTH*i+j];

			Memory[256*16+BUS_WIDTH*i+j]	=	INIT_10[BUS_WIDTH*i+j];
			Memory[256*17+BUS_WIDTH*i+j]	=	INIT_11[BUS_WIDTH*i+j];
			Memory[256*18+BUS_WIDTH*i+j]	=	INIT_12[BUS_WIDTH*i+j];
			Memory[256*19+BUS_WIDTH*i+j]	=	INIT_13[BUS_WIDTH*i+j];
			Memory[256*20+BUS_WIDTH*i+j]	=	INIT_14[BUS_WIDTH*i+j];
			Memory[256*21+BUS_WIDTH*i+j]	=	INIT_15[BUS_WIDTH*i+j];
			Memory[256*22+BUS_WIDTH*i+j]	=	INIT_16[BUS_WIDTH*i+j];
			Memory[256*23+BUS_WIDTH*i+j]	=	INIT_17[BUS_WIDTH*i+j];
			Memory[256*24+BUS_WIDTH*i+j]	=	INIT_18[BUS_WIDTH*i+j];
			Memory[256*25+BUS_WIDTH*i+j]	=	INIT_19[BUS_WIDTH*i+j];
			Memory[256*26+BUS_WIDTH*i+j]	=	INIT_1A[BUS_WIDTH*i+j];
			Memory[256*27+BUS_WIDTH*i+j]	=	INIT_1B[BUS_WIDTH*i+j];
			Memory[256*28+BUS_WIDTH*i+j]	=	INIT_1C[BUS_WIDTH*i+j];
			Memory[256*29+BUS_WIDTH*i+j]	=	INIT_1D[BUS_WIDTH*i+j];
			Memory[256*30+BUS_WIDTH*i+j]	=	INIT_1E[BUS_WIDTH*i+j];
			Memory[256*31+BUS_WIDTH*i+j]	=	INIT_1F[BUS_WIDTH*i+j];

			Memory[256*32+BUS_WIDTH*i+j]	=	INIT_20[BUS_WIDTH*i+j];
			Memory[256*33+BUS_WIDTH*i+j]	=	INIT_21[BUS_WIDTH*i+j];
			Memory[256*34+BUS_WIDTH*i+j]	=	INIT_22[BUS_WIDTH*i+j];
			Memory[256*35+BUS_WIDTH*i+j]	=	INIT_23[BUS_WIDTH*i+j];
			Memory[256*36+BUS_WIDTH*i+j]	=	INIT_24[BUS_WIDTH*i+j];
			Memory[256*37+BUS_WIDTH*i+j]	=	INIT_25[BUS_WIDTH*i+j];
			Memory[256*38+BUS_WIDTH*i+j]	=	INIT_26[BUS_WIDTH*i+j];
			Memory[256*39+BUS_WIDTH*i+j]	=	INIT_27[BUS_WIDTH*i+j];
			Memory[256*40+BUS_WIDTH*i+j]	=	INIT_28[BUS_WIDTH*i+j];
			Memory[256*41+BUS_WIDTH*i+j]	=	INIT_29[BUS_WIDTH*i+j];
			Memory[256*42+BUS_WIDTH*i+j]	=	INIT_2A[BUS_WIDTH*i+j];
			Memory[256*43+BUS_WIDTH*i+j]	=	INIT_2B[BUS_WIDTH*i+j];
			Memory[256*44+BUS_WIDTH*i+j]	=	INIT_2C[BUS_WIDTH*i+j];
			Memory[256*45+BUS_WIDTH*i+j]	=	INIT_2D[BUS_WIDTH*i+j];
			Memory[256*46+BUS_WIDTH*i+j]	=	INIT_2E[BUS_WIDTH*i+j];
			Memory[256*47+BUS_WIDTH*i+j]	=	INIT_2F[BUS_WIDTH*i+j];

			Memory[256*48+BUS_WIDTH*i+j]	=	INIT_30[BUS_WIDTH*i+j];
			Memory[256*49+BUS_WIDTH*i+j]	=	INIT_31[BUS_WIDTH*i+j];
			Memory[256*50+BUS_WIDTH*i+j]	=	INIT_32[BUS_WIDTH*i+j];
			Memory[256*51+BUS_WIDTH*i+j]	=	INIT_33[BUS_WIDTH*i+j];
			Memory[256*52+BUS_WIDTH*i+j]	=	INIT_34[BUS_WIDTH*i+j];
			Memory[256*53+BUS_WIDTH*i+j]	=	INIT_35[BUS_WIDTH*i+j];
			Memory[256*54+BUS_WIDTH*i+j]	=	INIT_36[BUS_WIDTH*i+j];
			Memory[256*55+BUS_WIDTH*i+j]	=	INIT_37[BUS_WIDTH*i+j];
			Memory[256*56+BUS_WIDTH*i+j]	=	INIT_38[BUS_WIDTH*i+j];
			Memory[256*57+BUS_WIDTH*i+j]	=	INIT_39[BUS_WIDTH*i+j];
			Memory[256*58+BUS_WIDTH*i+j]	=	INIT_3A[BUS_WIDTH*i+j];
			Memory[256*59+BUS_WIDTH*i+j]	=	INIT_3B[BUS_WIDTH*i+j];
			Memory[256*60+BUS_WIDTH*i+j]	=	INIT_3C[BUS_WIDTH*i+j];
			Memory[256*61+BUS_WIDTH*i+j]	=	INIT_3D[BUS_WIDTH*i+j];
			Memory[256*62+BUS_WIDTH*i+j]	=	INIT_3E[BUS_WIDTH*i+j];
			Memory[256*63+BUS_WIDTH*i+j]	=	INIT_3F[BUS_WIDTH*i+j];

		end 
	end

end

assign Address_Collision_Detected = ((RE & WE & WCLKE & RCLKE)&(WADDR == RADDR)); 

always @(WCLK or WCLKE) 
begin 
	if(~WCLK)
	WCLKE_sync = WCLKE;   	
end 

always @(RCLK or RCLKE) 
begin 
	if (~RCLK)
	RCLKE_sync = RCLKE; 	
end 

assign WCLK_g = WCLK & WCLKE_sync;
assign RCLK_g = RCLK & RCLKE_sync;


always @(posedge WCLK_g) begin
	time_WCLK = $time;
end

always @(posedge RCLK_g) begin
    	time_RCLK = $time;
end
integer	SB_RAM1024x16_RDATA_log_file;					//.....................
initial	SB_RAM1024x16_RDATA_log_file=("SB_RAM1024x16_RDATA_log_file.txt");	//.....................
always @(posedge WCLK_g) begin

	Time_Collision_Detected = Check_Timed_Window_Violation(time_WCLK,time_RCLK,COLLISION_TIME_WINDOW);
        if (Time_Collision_Detected & Address_Collision_Detected)begin
        	$display("Warning: Write-Read collision detected, Data read value is XXXX\n");
 		$display("WCLK Time: %.3f   RCLK Time:%.3f  ",time_WCLK, time_RCLK,"WADDR: %d   RADDR:%d\n",WADDR, RADDR); 
 		$fdisplay(SB_RAM1024x16_RDATA_log_file,"Warning: Write-Read collision detected, Data read value is XXXX\n");
		$fdisplay(SB_RAM1024x16_RDATA_log_file,"WCLK Time: %.3f   RCLK Time:%.3f  ",time_WCLK, time_RCLK, "WADDR: %d   RADDR:%d\n",WADDR, RADDR); 	
 		-> Collision_e;
	end
end

//	code modify for universal verilog compiler

always @ (posedge WCLK_g)
begin
	if	(WE)
	begin
		-> Write_e;
		for	(i=0;i<=BUS_WIDTH-1; i=i+1)
		begin
			if	(MASK[i] !=1)
				Memory[WADDR*BUS_WIDTH+i]	<=	WDATA[i];
			else
				Memory[WADDR*BUS_WIDTH+i]	<=	Memory[WADDR*BUS_WIDTH+i];
		end
	end
end

reg	[15:0]	RDATA = 0;

// Look at the rising edge of the clock

always @ (posedge RCLK_g)
begin
	if	(RE)
	begin
		-> Read_e;
		if	(Time_Collision_Detected & Address_Collision_Detected) 
			RDATA <= 16'hXXXX;
		else
			for	(i=0;i<=BUS_WIDTH-1;i=i+1)
				RDATA[i]	<= Memory[RADDR*BUS_WIDTH+i];
	end
end

`ifdef TIMINGCHECK
specify
   (RCLK *> RDATA[0]) = (1.0, 1.0);
   (RCLK *> RDATA[1]) = (1.0, 1.0);
   (RCLK *> RDATA[2]) = (1.0, 1.0);
   (RCLK *> RDATA[3]) = (1.0, 1.0);
   (RCLK *> RDATA[4]) = (1.0, 1.0);
   (RCLK *> RDATA[5]) = (1.0, 1.0);
   (RCLK *> RDATA[6]) = (1.0, 1.0);
   (RCLK *> RDATA[7]) = (1.0, 1.0);
   (RCLK *> RDATA[8]) = (1.0, 1.0);
   (RCLK *> RDATA[9]) = (1.0, 1.0);
   (RCLK *> RDATA[10]) = (1.0, 1.0);
   (RCLK *> RDATA[11]) = (1.0, 1.0);
   (RCLK *> RDATA[12]) = (1.0, 1.0);
   (RCLK *> RDATA[13]) = (1.0, 1.0);
   (RCLK *> RDATA[14]) = (1.0, 1.0);
   (RCLK *> RDATA[15]) = (1.0, 1.0);
   $setup(posedge MASK[0], posedge WCLK, 1.0);
   $setup(negedge MASK[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[0], 1.0);
   $hold(posedge WCLK, negedge MASK[0], 1.0);
   $setup(posedge MASK[1], posedge WCLK, 1.0);
   $setup(negedge MASK[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[1], 1.0);
   $hold(posedge WCLK, negedge MASK[1], 1.0);
   $setup(posedge MASK[2], posedge WCLK, 1.0);
   $setup(negedge MASK[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[2], 1.0);
   $hold(posedge WCLK, negedge MASK[2], 1.0);
   $setup(posedge MASK[3], posedge WCLK, 1.0);
   $setup(negedge MASK[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[3], 1.0);
   $hold(posedge WCLK, negedge MASK[3], 1.0);
   $setup(posedge MASK[4], posedge WCLK, 1.0);
   $setup(negedge MASK[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[4], 1.0);
   $hold(posedge WCLK, negedge MASK[4], 1.0);
   $setup(posedge MASK[5], posedge WCLK, 1.0);
   $setup(negedge MASK[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[5], 1.0);
   $hold(posedge WCLK, negedge MASK[5], 1.0);
   $setup(posedge MASK[6], posedge WCLK, 1.0);
   $setup(negedge MASK[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[6], 1.0);
   $hold(posedge WCLK, negedge MASK[6], 1.0);
   $setup(posedge MASK[7], posedge WCLK, 1.0);
   $setup(negedge MASK[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[7], 1.0);
   $hold(posedge WCLK, negedge MASK[7], 1.0);
   $setup(posedge MASK[8], posedge WCLK, 1.0);
   $setup(negedge MASK[8], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[8], 1.0);
   $hold(posedge WCLK, negedge MASK[8], 1.0);
   $setup(posedge MASK[9], posedge WCLK, 1.0);
   $setup(negedge MASK[9], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[9], 1.0);
   $hold(posedge WCLK, negedge MASK[9], 1.0);
   $setup(posedge MASK[10], posedge WCLK, 1.0);
   $setup(negedge MASK[10], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[10], 1.0);
   $hold(posedge WCLK, negedge MASK[10], 1.0);
   $setup(posedge MASK[11], posedge WCLK, 1.0);
   $setup(negedge MASK[11], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[11], 1.0);
   $hold(posedge WCLK, negedge MASK[11], 1.0);
   $setup(posedge MASK[12], posedge WCLK, 1.0);
   $setup(negedge MASK[12], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[12], 1.0);
   $hold(posedge WCLK, negedge MASK[12], 1.0);
   $setup(posedge MASK[13], posedge WCLK, 1.0);
   $setup(negedge MASK[13], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[13], 1.0);
   $hold(posedge WCLK, negedge MASK[13], 1.0);
   $setup(posedge MASK[14], posedge WCLK, 1.0);
   $setup(negedge MASK[14], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[14], 1.0);
   $hold(posedge WCLK, negedge MASK[14], 1.0);
   $setup(posedge MASK[15], posedge WCLK, 1.0);
   $setup(negedge MASK[15], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[15], 1.0);
   $hold(posedge WCLK, negedge MASK[15], 1.0);
   $setup(posedge WADDR[0], posedge WCLK, 1.0);
   $setup(negedge WADDR[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[0], 1.0);
   $hold(posedge WCLK, negedge WADDR[0], 1.0);
   $setup(posedge WADDR[1], posedge WCLK, 1.0);
   $setup(negedge WADDR[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[1], 1.0);
   $hold(posedge WCLK, negedge WADDR[1], 1.0);
   $setup(posedge WADDR[2], posedge WCLK, 1.0);
   $setup(negedge WADDR[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[2], 1.0);
   $hold(posedge WCLK, negedge WADDR[2], 1.0);
   $setup(posedge WADDR[3], posedge WCLK, 1.0);
   $setup(negedge WADDR[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[3], 1.0);
   $hold(posedge WCLK, negedge WADDR[3], 1.0);
   $setup(posedge WADDR[4], posedge WCLK, 1.0);
   $setup(negedge WADDR[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[4], 1.0);
   $hold(posedge WCLK, negedge WADDR[4], 1.0);
   $setup(posedge WADDR[5], posedge WCLK, 1.0);
   $setup(negedge WADDR[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[5], 1.0);
   $hold(posedge WCLK, negedge WADDR[5], 1.0);
   $setup(posedge WADDR[6], posedge WCLK, 1.0);
   $setup(negedge WADDR[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[6], 1.0);
   $hold(posedge WCLK, negedge WADDR[6], 1.0);
   $setup(posedge WADDR[7], posedge WCLK, 1.0);
   $setup(negedge WADDR[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[7], 1.0);
   $hold(posedge WCLK, negedge WADDR[7], 1.0);
   $setup(posedge WADDR[8], posedge WCLK, 1.0);
   $setup(negedge WADDR[8], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[8], 1.0);
   $hold(posedge WCLK, negedge WADDR[8], 1.0);
   $setup(posedge WADDR[9], posedge WCLK, 1.0);
   $setup(negedge WADDR[9], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[9], 1.0);
   $hold(posedge WCLK, negedge WADDR[9], 1.0);
   $setup(posedge WDATA[0], posedge WCLK, 1.0);
   $setup(negedge WDATA[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[0], 1.0);
   $hold(posedge WCLK, negedge WDATA[0], 1.0);
   $setup(posedge WDATA[1], posedge WCLK, 1.0);
   $setup(negedge WDATA[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[1], 1.0);
   $hold(posedge WCLK, negedge WDATA[1], 1.0);
   $setup(posedge WDATA[2], posedge WCLK, 1.0);
   $setup(negedge WDATA[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[2], 1.0);
   $hold(posedge WCLK, negedge WDATA[2], 1.0);
   $setup(posedge WDATA[3], posedge WCLK, 1.0);
   $setup(negedge WDATA[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[3], 1.0);
   $hold(posedge WCLK, negedge WDATA[3], 1.0);
   $setup(posedge WDATA[4], posedge WCLK, 1.0);
   $setup(negedge WDATA[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[4], 1.0);
   $hold(posedge WCLK, negedge WDATA[4], 1.0);
   $setup(posedge WDATA[5], posedge WCLK, 1.0);
   $setup(negedge WDATA[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[5], 1.0);
   $hold(posedge WCLK, negedge WDATA[5], 1.0);
   $setup(posedge WDATA[6], posedge WCLK, 1.0);
   $setup(negedge WDATA[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[6], 1.0);
   $hold(posedge WCLK, negedge WDATA[6], 1.0);
   $setup(posedge WDATA[7], posedge WCLK, 1.0);
   $setup(negedge WDATA[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[7], 1.0);
   $hold(posedge WCLK, negedge WDATA[7], 1.0);
   $setup(posedge WDATA[8], posedge WCLK, 1.0);
   $setup(negedge WDATA[8], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[8], 1.0);
   $hold(posedge WCLK, negedge WDATA[8], 1.0);
   $setup(posedge WDATA[9], posedge WCLK, 1.0);
   $setup(negedge WDATA[9], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[9], 1.0);
   $hold(posedge WCLK, negedge WDATA[9], 1.0);
   $setup(posedge WDATA[10], posedge WCLK, 1.0);
   $setup(negedge WDATA[10], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[10], 1.0);
   $hold(posedge WCLK, negedge WDATA[10], 1.0);
   $setup(posedge WDATA[11], posedge WCLK, 1.0);
   $setup(negedge WDATA[11], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[11], 1.0);
   $hold(posedge WCLK, negedge WDATA[11], 1.0);
   $setup(posedge WDATA[12], posedge WCLK, 1.0);
   $setup(negedge WDATA[12], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[12], 1.0);
   $hold(posedge WCLK, negedge WDATA[12], 1.0);
   $setup(posedge WDATA[13], posedge WCLK, 1.0);
   $setup(negedge WDATA[13], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[13], 1.0);
   $hold(posedge WCLK, negedge WDATA[13], 1.0);
   $setup(posedge WDATA[14], posedge WCLK, 1.0);
   $setup(negedge WDATA[14], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[14], 1.0);
   $hold(posedge WCLK, negedge WDATA[14], 1.0);
   $setup(posedge WDATA[15], posedge WCLK, 1.0);
   $setup(negedge WDATA[15], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[15], 1.0);
   $hold(posedge WCLK, negedge WDATA[15], 1.0);
   $setup(posedge WCLKE, posedge WCLK, 1.0);
   $setup(negedge WCLKE, posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WCLKE, 1.0);
   $hold(posedge WCLK, negedge WCLKE, 1.0);
   $setup(posedge WE, posedge WCLK, 1.0);
   $setup(negedge WE, posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WE, 1.0);
   $hold(posedge WCLK, negedge WE, 1.0);
   $setup(posedge RADDR[0], posedge RCLK, 1.0);
   $setup(negedge RADDR[0], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[0], 1.0);
   $hold(posedge RCLK, negedge RADDR[0], 1.0);
   $setup(posedge RADDR[1], posedge RCLK, 1.0);
   $setup(negedge RADDR[1], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[1], 1.0);
   $hold(posedge RCLK, negedge RADDR[1], 1.0);
   $setup(posedge RADDR[2], posedge RCLK, 1.0);
   $setup(negedge RADDR[2], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[2], 1.0);
   $hold(posedge RCLK, negedge RADDR[2], 1.0);
   $setup(posedge RADDR[3], posedge RCLK, 1.0);
   $setup(negedge RADDR[3], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[3], 1.0);
   $hold(posedge RCLK, negedge RADDR[3], 1.0);
   $setup(posedge RADDR[4], posedge RCLK, 1.0);
   $setup(negedge RADDR[4], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[4], 1.0);
   $hold(posedge RCLK, negedge RADDR[4], 1.0);
   $setup(posedge RADDR[5], posedge RCLK, 1.0);
   $setup(negedge RADDR[5], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[5], 1.0);
   $hold(posedge RCLK, negedge RADDR[5], 1.0);
   $setup(posedge RADDR[6], posedge RCLK, 1.0);
   $setup(negedge RADDR[6], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[6], 1.0);
   $hold(posedge RCLK, negedge RADDR[6], 1.0);
   $setup(posedge RADDR[7], posedge RCLK, 1.0);
   $setup(negedge RADDR[7], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[7], 1.0);
   $hold(posedge RCLK, negedge RADDR[7], 1.0);
   $setup(posedge RADDR[8], posedge RCLK, 1.0);
   $setup(negedge RADDR[8], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[8], 1.0);
   $hold(posedge RCLK, negedge RADDR[8], 1.0);
   $setup(posedge RADDR[9], posedge RCLK, 1.0);
   $setup(negedge RADDR[9], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[9], 1.0);
   $hold(posedge RCLK, negedge RADDR[9], 1.0);
   $setup(posedge RCLKE, posedge RCLK, 1.0);
   $setup(negedge RCLKE, posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RCLKE, 1.0);
   $hold(posedge RCLK, negedge RCLKE, 1.0);
   $setup(posedge RE, posedge RCLK, 1.0);
   $setup(negedge RE, posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RE, 1.0);
   $hold(posedge RCLK, negedge RE, 1.0);
endspecify
`endif

endmodule   //SB_RAM1024x16     
  
//---------------------------------------
// 	--- SB_RAM1024x16NR
//---------------------------------------
`timescale 1ps/1ps
module SB_RAM1024x16NR ( RDATA, RCLKN, RCLKE, RE, RADDR, WCLK, WCLKE, WE, WADDR, MASK, WDATA );  

output	[15:0]	RDATA;  
input         	RCLKN;   
input           RCLKE; 
input           RE; 
input	[9:0]   RADDR; 
input           WCLK; 
input           WCLKE; 
input           WE; 
input 	[9:0]   WADDR; 
input	[15:0]	MASK; 
input 	[15:0]	WDATA; 


parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

wire RCLK;
assign (weak0, weak1) RCLKE =1'b1 ;
assign (weak0, weak1) RE =1'b0 ;
assign (weak0, weak1) WCLKE =1'b1 ;
assign (weak0, weak1) WE =1'b0 ;
assign RCLK = ~RCLKN;

SB_RAM1024x16 sb_ram1024x16r_inst (
	.RDATA(RDATA),
	.RCLK(RCLK),
	.RCLKE(RCLKE),
	.RE(RE),
	.RADDR(RADDR),
	.WCLK(WCLK),
	.WCLKE(WCLKE),
	.WE(WE),
	.WADDR(WADDR),
	.MASK(MASK),
	.WDATA(WDATA));

defparam sb_ram1024x16r_inst.INIT_0 = INIT_0;
defparam sb_ram1024x16r_inst.INIT_1 = INIT_1;
defparam sb_ram1024x16r_inst.INIT_2 = INIT_2;
defparam sb_ram1024x16r_inst.INIT_3 = INIT_3;
defparam sb_ram1024x16r_inst.INIT_4 = INIT_4;
defparam sb_ram1024x16r_inst.INIT_5 = INIT_5;
defparam sb_ram1024x16r_inst.INIT_6 = INIT_6;
defparam sb_ram1024x16r_inst.INIT_7 = INIT_7;
defparam sb_ram1024x16r_inst.INIT_8 = INIT_8;
defparam sb_ram1024x16r_inst.INIT_9 = INIT_9;
defparam sb_ram1024x16r_inst.INIT_A = INIT_A;
defparam sb_ram1024x16r_inst.INIT_B = INIT_B;
defparam sb_ram1024x16r_inst.INIT_C = INIT_C;
defparam sb_ram1024x16r_inst.INIT_D = INIT_D;
defparam sb_ram1024x16r_inst.INIT_E = INIT_E;
defparam sb_ram1024x16r_inst.INIT_F = INIT_F;

defparam sb_ram1024x16r_inst.INIT_10 = INIT_10;
defparam sb_ram1024x16r_inst.INIT_11 = INIT_11;
defparam sb_ram1024x16r_inst.INIT_12 = INIT_12;
defparam sb_ram1024x16r_inst.INIT_13 = INIT_13;
defparam sb_ram1024x16r_inst.INIT_14 = INIT_14;
defparam sb_ram1024x16r_inst.INIT_15 = INIT_15;
defparam sb_ram1024x16r_inst.INIT_16 = INIT_16;
defparam sb_ram1024x16r_inst.INIT_17 = INIT_17;
defparam sb_ram1024x16r_inst.INIT_18 = INIT_18;
defparam sb_ram1024x16r_inst.INIT_19 = INIT_19;
defparam sb_ram1024x16r_inst.INIT_1A = INIT_1A;
defparam sb_ram1024x16r_inst.INIT_1B = INIT_1B;
defparam sb_ram1024x16r_inst.INIT_1C = INIT_1C;
defparam sb_ram1024x16r_inst.INIT_1D = INIT_1D;
defparam sb_ram1024x16r_inst.INIT_1E = INIT_1E;
defparam sb_ram1024x16r_inst.INIT_1F = INIT_1F;

defparam sb_ram1024x16r_inst.INIT_20 = INIT_20;
defparam sb_ram1024x16r_inst.INIT_21 = INIT_21;
defparam sb_ram1024x16r_inst.INIT_22 = INIT_22;
defparam sb_ram1024x16r_inst.INIT_23 = INIT_23;
defparam sb_ram1024x16r_inst.INIT_24 = INIT_24;
defparam sb_ram1024x16r_inst.INIT_25 = INIT_25;
defparam sb_ram1024x16r_inst.INIT_26 = INIT_26;
defparam sb_ram1024x16r_inst.INIT_27 = INIT_27;
defparam sb_ram1024x16r_inst.INIT_28 = INIT_28;
defparam sb_ram1024x16r_inst.INIT_29 = INIT_29;
defparam sb_ram1024x16r_inst.INIT_2A = INIT_2A;
defparam sb_ram1024x16r_inst.INIT_2B = INIT_2B;
defparam sb_ram1024x16r_inst.INIT_2C = INIT_2C;
defparam sb_ram1024x16r_inst.INIT_2D = INIT_2D;
defparam sb_ram1024x16r_inst.INIT_2E = INIT_2E;
defparam sb_ram1024x16r_inst.INIT_2F = INIT_2F;

defparam sb_ram1024x16r_inst.INIT_30 = INIT_30;
defparam sb_ram1024x16r_inst.INIT_31 = INIT_31;
defparam sb_ram1024x16r_inst.INIT_32 = INIT_32;
defparam sb_ram1024x16r_inst.INIT_33 = INIT_33;
defparam sb_ram1024x16r_inst.INIT_34 = INIT_34;
defparam sb_ram1024x16r_inst.INIT_35 = INIT_35;
defparam sb_ram1024x16r_inst.INIT_36 = INIT_36;
defparam sb_ram1024x16r_inst.INIT_37 = INIT_37;
defparam sb_ram1024x16r_inst.INIT_38 = INIT_38;
defparam sb_ram1024x16r_inst.INIT_39 = INIT_39;
defparam sb_ram1024x16r_inst.INIT_3A = INIT_3A;
defparam sb_ram1024x16r_inst.INIT_3B = INIT_3B;
defparam sb_ram1024x16r_inst.INIT_3C = INIT_3C;
defparam sb_ram1024x16r_inst.INIT_3D = INIT_3D;
defparam sb_ram1024x16r_inst.INIT_3E = INIT_3E;
defparam sb_ram1024x16r_inst.INIT_3F = INIT_3F;


`ifdef TIMINGCHECK
specify
   (RCLKN *> RDATA[0]) = (1.0, 1.0);
   (RCLKN *> RDATA[1]) = (1.0, 1.0);
   (RCLKN *> RDATA[2]) = (1.0, 1.0);
   (RCLKN *> RDATA[3]) = (1.0, 1.0);
   (RCLKN *> RDATA[4]) = (1.0, 1.0);
   (RCLKN *> RDATA[5]) = (1.0, 1.0);
   (RCLKN *> RDATA[6]) = (1.0, 1.0);
   (RCLKN *> RDATA[7]) = (1.0, 1.0);
   (RCLKN *> RDATA[8]) = (1.0, 1.0);
   (RCLKN *> RDATA[9]) = (1.0, 1.0);
   (RCLKN *> RDATA[10]) = (1.0, 1.0);
   (RCLKN *> RDATA[11]) = (1.0, 1.0);
   (RCLKN *> RDATA[12]) = (1.0, 1.0);
   (RCLKN *> RDATA[13]) = (1.0, 1.0);
   (RCLKN *> RDATA[14]) = (1.0, 1.0);
   (RCLKN *> RDATA[15]) = (1.0, 1.0);
   $setup(posedge MASK[0], posedge WCLK, 1.0);
   $setup(negedge MASK[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[0], 1.0);
   $hold(posedge WCLK, negedge MASK[0], 1.0);
   $setup(posedge MASK[1], posedge WCLK, 1.0);
   $setup(negedge MASK[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[1], 1.0);
   $hold(posedge WCLK, negedge MASK[1], 1.0);
   $setup(posedge MASK[2], posedge WCLK, 1.0);
   $setup(negedge MASK[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[2], 1.0);
   $hold(posedge WCLK, negedge MASK[2], 1.0);
   $setup(posedge MASK[3], posedge WCLK, 1.0);
   $setup(negedge MASK[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[3], 1.0);
   $hold(posedge WCLK, negedge MASK[3], 1.0);
   $setup(posedge MASK[4], posedge WCLK, 1.0);
   $setup(negedge MASK[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[4], 1.0);
   $hold(posedge WCLK, negedge MASK[4], 1.0);
   $setup(posedge MASK[5], posedge WCLK, 1.0);
   $setup(negedge MASK[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[5], 1.0);
   $hold(posedge WCLK, negedge MASK[5], 1.0);
   $setup(posedge MASK[6], posedge WCLK, 1.0);
   $setup(negedge MASK[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[6], 1.0);
   $hold(posedge WCLK, negedge MASK[6], 1.0);
   $setup(posedge MASK[7], posedge WCLK, 1.0);
   $setup(negedge MASK[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[7], 1.0);
   $hold(posedge WCLK, negedge MASK[7], 1.0);
   $setup(posedge MASK[8], posedge WCLK, 1.0);
   $setup(negedge MASK[8], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[8], 1.0);
   $hold(posedge WCLK, negedge MASK[8], 1.0);
   $setup(posedge MASK[9], posedge WCLK, 1.0);
   $setup(negedge MASK[9], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[9], 1.0);
   $hold(posedge WCLK, negedge MASK[9], 1.0);
   $setup(posedge MASK[10], posedge WCLK, 1.0);
   $setup(negedge MASK[10], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[10], 1.0);
   $hold(posedge WCLK, negedge MASK[10], 1.0);
   $setup(posedge MASK[11], posedge WCLK, 1.0);
   $setup(negedge MASK[11], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[11], 1.0);
   $hold(posedge WCLK, negedge MASK[11], 1.0);
   $setup(posedge MASK[12], posedge WCLK, 1.0);
   $setup(negedge MASK[12], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[12], 1.0);
   $hold(posedge WCLK, negedge MASK[12], 1.0);
   $setup(posedge MASK[13], posedge WCLK, 1.0);
   $setup(negedge MASK[13], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[13], 1.0);
   $hold(posedge WCLK, negedge MASK[13], 1.0);
   $setup(posedge MASK[14], posedge WCLK, 1.0);
   $setup(negedge MASK[14], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[14], 1.0);
   $hold(posedge WCLK, negedge MASK[14], 1.0);
   $setup(posedge MASK[15], posedge WCLK, 1.0);
   $setup(negedge MASK[15], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[15], 1.0);
   $hold(posedge WCLK, negedge MASK[15], 1.0);
   $setup(posedge WADDR[0], posedge WCLK, 1.0);
   $setup(negedge WADDR[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[0], 1.0);
   $hold(posedge WCLK, negedge WADDR[0], 1.0);
   $setup(posedge WADDR[1], posedge WCLK, 1.0);
   $setup(negedge WADDR[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[1], 1.0);
   $hold(posedge WCLK, negedge WADDR[1], 1.0);
   $setup(posedge WADDR[2], posedge WCLK, 1.0);
   $setup(negedge WADDR[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[2], 1.0);
   $hold(posedge WCLK, negedge WADDR[2], 1.0);
   $setup(posedge WADDR[3], posedge WCLK, 1.0);
   $setup(negedge WADDR[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[3], 1.0);
   $hold(posedge WCLK, negedge WADDR[3], 1.0);
   $setup(posedge WADDR[4], posedge WCLK, 1.0);
   $setup(negedge WADDR[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[4], 1.0);
   $hold(posedge WCLK, negedge WADDR[4], 1.0);
   $setup(posedge WADDR[5], posedge WCLK, 1.0);
   $setup(negedge WADDR[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[5], 1.0);
   $hold(posedge WCLK, negedge WADDR[5], 1.0);
   $setup(posedge WADDR[6], posedge WCLK, 1.0);
   $setup(negedge WADDR[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[6], 1.0);
   $hold(posedge WCLK, negedge WADDR[6], 1.0);
   $setup(posedge WADDR[7], posedge WCLK, 1.0);
   $setup(negedge WADDR[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[7], 1.0);
   $hold(posedge WCLK, negedge WADDR[7], 1.0);
   $setup(posedge WADDR[8], posedge WCLK, 1.0);
   $setup(negedge WADDR[8], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[8], 1.0);
   $hold(posedge WCLK, negedge WADDR[8], 1.0);
   $setup(posedge WADDR[9], posedge WCLK, 1.0);
   $setup(negedge WADDR[9], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[9], 1.0);
   $hold(posedge WCLK, negedge WADDR[9], 1.0);
   $setup(posedge WDATA[0], posedge WCLK, 1.0);
   $setup(negedge WDATA[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[0], 1.0);
   $hold(posedge WCLK, negedge WDATA[0], 1.0);
   $setup(posedge WDATA[1], posedge WCLK, 1.0);
   $setup(negedge WDATA[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[1], 1.0);
   $hold(posedge WCLK, negedge WDATA[1], 1.0);
   $setup(posedge WDATA[2], posedge WCLK, 1.0);
   $setup(negedge WDATA[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[2], 1.0);
   $hold(posedge WCLK, negedge WDATA[2], 1.0);
   $setup(posedge WDATA[3], posedge WCLK, 1.0);
   $setup(negedge WDATA[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[3], 1.0);
   $hold(posedge WCLK, negedge WDATA[3], 1.0);
   $setup(posedge WDATA[4], posedge WCLK, 1.0);
   $setup(negedge WDATA[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[4], 1.0);
   $hold(posedge WCLK, negedge WDATA[4], 1.0);
   $setup(posedge WDATA[5], posedge WCLK, 1.0);
   $setup(negedge WDATA[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[5], 1.0);
   $hold(posedge WCLK, negedge WDATA[5], 1.0);
   $setup(posedge WDATA[6], posedge WCLK, 1.0);
   $setup(negedge WDATA[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[6], 1.0);
   $hold(posedge WCLK, negedge WDATA[6], 1.0);
   $setup(posedge WDATA[7], posedge WCLK, 1.0);
   $setup(negedge WDATA[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[7], 1.0);
   $hold(posedge WCLK, negedge WDATA[7], 1.0);
   $setup(posedge WDATA[8], posedge WCLK, 1.0);
   $setup(negedge WDATA[8], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[8], 1.0);
   $hold(posedge WCLK, negedge WDATA[8], 1.0);
   $setup(posedge WDATA[9], posedge WCLK, 1.0);
   $setup(negedge WDATA[9], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[9], 1.0);
   $hold(posedge WCLK, negedge WDATA[9], 1.0);
   $setup(posedge WDATA[10], posedge WCLK, 1.0);
   $setup(negedge WDATA[10], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[10], 1.0);
   $hold(posedge WCLK, negedge WDATA[10], 1.0);
   $setup(posedge WDATA[11], posedge WCLK, 1.0);
   $setup(negedge WDATA[11], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[11], 1.0);
   $hold(posedge WCLK, negedge WDATA[11], 1.0);
   $setup(posedge WDATA[12], posedge WCLK, 1.0);
   $setup(negedge WDATA[12], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[12], 1.0);
   $hold(posedge WCLK, negedge WDATA[12], 1.0);
   $setup(posedge WDATA[13], posedge WCLK, 1.0);
   $setup(negedge WDATA[13], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[13], 1.0);
   $hold(posedge WCLK, negedge WDATA[13], 1.0);
   $setup(posedge WDATA[14], posedge WCLK, 1.0);
   $setup(negedge WDATA[14], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[14], 1.0);
   $hold(posedge WCLK, negedge WDATA[14], 1.0);
   $setup(posedge WDATA[15], posedge WCLK, 1.0);
   $setup(negedge WDATA[15], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[15], 1.0);
   $hold(posedge WCLK, negedge WDATA[15], 1.0);
   $setup(posedge WCLKE, posedge WCLK, 1.0);
   $setup(negedge WCLKE, posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WCLKE, 1.0);
   $hold(posedge WCLK, negedge WCLKE, 1.0);
   $setup(posedge WE, posedge WCLK, 1.0);
   $setup(negedge WE, posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WE, 1.0);
   $hold(posedge WCLK, negedge WE, 1.0);
   $setup(posedge RADDR[0], posedge RCLKN, 1.0);
   $setup(negedge RADDR[0], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[0], 1.0);
   $hold(posedge RCLKN, negedge RADDR[0], 1.0);
   $setup(posedge RADDR[1], posedge RCLKN, 1.0);
   $setup(negedge RADDR[1], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[1], 1.0);
   $hold(posedge RCLKN, negedge RADDR[1], 1.0);
   $setup(posedge RADDR[2], posedge RCLKN, 1.0);
   $setup(negedge RADDR[2], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[2], 1.0);
   $hold(posedge RCLKN, negedge RADDR[2], 1.0);
   $setup(posedge RADDR[3], posedge RCLKN, 1.0);
   $setup(negedge RADDR[3], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[3], 1.0);
   $hold(posedge RCLKN, negedge RADDR[3], 1.0);
   $setup(posedge RADDR[4], posedge RCLKN, 1.0);
   $setup(negedge RADDR[4], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[4], 1.0);
   $hold(posedge RCLKN, negedge RADDR[4], 1.0);
   $setup(posedge RADDR[5], posedge RCLKN, 1.0);
   $setup(negedge RADDR[5], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[5], 1.0);
   $hold(posedge RCLKN, negedge RADDR[5], 1.0);
   $setup(posedge RADDR[6], posedge RCLKN, 1.0);
   $setup(negedge RADDR[6], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[6], 1.0);
   $hold(posedge RCLKN, negedge RADDR[6], 1.0);
   $setup(posedge RADDR[7], posedge RCLKN, 1.0);
   $setup(negedge RADDR[7], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[7], 1.0);
   $hold(posedge RCLKN, negedge RADDR[7], 1.0);
   $setup(posedge RADDR[8], posedge RCLKN, 1.0);
   $setup(negedge RADDR[8], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[8], 1.0);
   $hold(posedge RCLKN, negedge RADDR[8], 1.0);
   $setup(posedge RADDR[9], posedge RCLKN, 1.0);
   $setup(negedge RADDR[9], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[9], 1.0);
   $hold(posedge RCLKN, negedge RADDR[9], 1.0);
   $setup(posedge RCLKE, posedge RCLKN, 1.0);
   $setup(negedge RCLKE, posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RCLKE, 1.0);
   $hold(posedge RCLKN, negedge RCLKE, 1.0);
   $setup(posedge RE, posedge RCLKN, 1.0);
   $setup(negedge RE, posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RE, 1.0);
   $hold(posedge RCLKN, negedge RE, 1.0);
endspecify
`endif

endmodule  //SB_RAM1024x16NR 

//---------------------------------------
//	--- SB_RAM1024x16NW
//---------------------------------------
`timescale 1ps/1ps
module SB_RAM1024x16NW  ( RDATA, RCLK, RCLKE, RE, RADDR, WCLKN, WCLKE, WE, WADDR, MASK, WDATA ); 

output	[15:0]	RDATA;  
input         	RCLK;   
input           RCLKE; 
input           RE; 
input	[9:0]   RADDR; 
input           WCLKN; 
input           WCLKE; 
input           WE; 
input 	[9:0]   WADDR; 
input	[15:0]	MASK; 
input 	[15:0]	WDATA; 
 
parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
 
wire WCLK;
assign (weak0, weak1) RCLKE =1'b1 ;
assign (weak0, weak1) RE =1'b0 ;
assign (weak0, weak1) WCLKE =1'b1 ;
assign (weak0, weak1) WE =1'b0 ;
assign WCLK = ~WCLKN;

SB_RAM1024x16 sb_ram1024x16w_inst (
	.RDATA(RDATA),
	.RCLK(RCLK),
	.RCLKE(RCLKE),
	.RE(RE),
	.RADDR(RADDR),
	.WCLK(WCLK),
	.WCLKE(WCLKE),
	.WE(WE),
	.WADDR(WADDR),
	.MASK(MASK),
	.WDATA(WDATA));

defparam sb_ram1024x16w_inst.INIT_0 = INIT_0;
defparam sb_ram1024x16w_inst.INIT_1 = INIT_1;
defparam sb_ram1024x16w_inst.INIT_2 = INIT_2;
defparam sb_ram1024x16w_inst.INIT_3 = INIT_3;
defparam sb_ram1024x16w_inst.INIT_4 = INIT_4;
defparam sb_ram1024x16w_inst.INIT_5 = INIT_5;
defparam sb_ram1024x16w_inst.INIT_6 = INIT_6;
defparam sb_ram1024x16w_inst.INIT_7 = INIT_7;
defparam sb_ram1024x16w_inst.INIT_8 = INIT_8;
defparam sb_ram1024x16w_inst.INIT_9 = INIT_9;
defparam sb_ram1024x16w_inst.INIT_A = INIT_A;
defparam sb_ram1024x16w_inst.INIT_B = INIT_B;
defparam sb_ram1024x16w_inst.INIT_C = INIT_C;
defparam sb_ram1024x16w_inst.INIT_D = INIT_D;
defparam sb_ram1024x16w_inst.INIT_E = INIT_E;
defparam sb_ram1024x16w_inst.INIT_F = INIT_F;

defparam sb_ram1024x16w_inst.INIT_10 = INIT_10;
defparam sb_ram1024x16w_inst.INIT_11 = INIT_11;
defparam sb_ram1024x16w_inst.INIT_12 = INIT_12;
defparam sb_ram1024x16w_inst.INIT_13 = INIT_13;
defparam sb_ram1024x16w_inst.INIT_14 = INIT_14;
defparam sb_ram1024x16w_inst.INIT_15 = INIT_15;
defparam sb_ram1024x16w_inst.INIT_16 = INIT_16;
defparam sb_ram1024x16w_inst.INIT_17 = INIT_17;
defparam sb_ram1024x16w_inst.INIT_18 = INIT_18;
defparam sb_ram1024x16w_inst.INIT_19 = INIT_19;
defparam sb_ram1024x16w_inst.INIT_1A = INIT_1A;
defparam sb_ram1024x16w_inst.INIT_1B = INIT_1B;
defparam sb_ram1024x16w_inst.INIT_1C = INIT_1C;
defparam sb_ram1024x16w_inst.INIT_1D = INIT_1D;
defparam sb_ram1024x16w_inst.INIT_1E = INIT_1E;
defparam sb_ram1024x16w_inst.INIT_1F = INIT_1F;

defparam sb_ram1024x16w_inst.INIT_20 = INIT_20;
defparam sb_ram1024x16w_inst.INIT_21 = INIT_21;
defparam sb_ram1024x16w_inst.INIT_22 = INIT_22;
defparam sb_ram1024x16w_inst.INIT_23 = INIT_23;
defparam sb_ram1024x16w_inst.INIT_24 = INIT_24;
defparam sb_ram1024x16w_inst.INIT_25 = INIT_25;
defparam sb_ram1024x16w_inst.INIT_26 = INIT_26;
defparam sb_ram1024x16w_inst.INIT_27 = INIT_27;
defparam sb_ram1024x16w_inst.INIT_28 = INIT_28;
defparam sb_ram1024x16w_inst.INIT_29 = INIT_29;
defparam sb_ram1024x16w_inst.INIT_2A = INIT_2A;
defparam sb_ram1024x16w_inst.INIT_2B = INIT_2B;
defparam sb_ram1024x16w_inst.INIT_2C = INIT_2C;
defparam sb_ram1024x16w_inst.INIT_2D = INIT_2D;
defparam sb_ram1024x16w_inst.INIT_2E = INIT_2E;
defparam sb_ram1024x16w_inst.INIT_2F = INIT_2F;

defparam sb_ram1024x16w_inst.INIT_30 = INIT_30;
defparam sb_ram1024x16w_inst.INIT_31 = INIT_31;
defparam sb_ram1024x16w_inst.INIT_32 = INIT_32;
defparam sb_ram1024x16w_inst.INIT_33 = INIT_33;
defparam sb_ram1024x16w_inst.INIT_34 = INIT_34;
defparam sb_ram1024x16w_inst.INIT_35 = INIT_35;
defparam sb_ram1024x16w_inst.INIT_36 = INIT_36;
defparam sb_ram1024x16w_inst.INIT_37 = INIT_37;
defparam sb_ram1024x16w_inst.INIT_38 = INIT_38;
defparam sb_ram1024x16w_inst.INIT_39 = INIT_39;
defparam sb_ram1024x16w_inst.INIT_3A = INIT_3A;
defparam sb_ram1024x16w_inst.INIT_3B = INIT_3B;
defparam sb_ram1024x16w_inst.INIT_3C = INIT_3C;
defparam sb_ram1024x16w_inst.INIT_3D = INIT_3D;
defparam sb_ram1024x16w_inst.INIT_3E = INIT_3E;
defparam sb_ram1024x16w_inst.INIT_3F = INIT_3F;

`ifdef TIMINGCHECK
specify
   (RCLK *> RDATA[0]) = (1.0, 1.0);
   (RCLK *> RDATA[1]) = (1.0, 1.0);
   (RCLK *> RDATA[2]) = (1.0, 1.0);
   (RCLK *> RDATA[3]) = (1.0, 1.0);
   (RCLK *> RDATA[4]) = (1.0, 1.0);
   (RCLK *> RDATA[5]) = (1.0, 1.0);
   (RCLK *> RDATA[6]) = (1.0, 1.0);
   (RCLK *> RDATA[7]) = (1.0, 1.0);
   (RCLK *> RDATA[8]) = (1.0, 1.0);
   (RCLK *> RDATA[9]) = (1.0, 1.0);
   (RCLK *> RDATA[10]) = (1.0, 1.0);
   (RCLK *> RDATA[11]) = (1.0, 1.0);
   (RCLK *> RDATA[12]) = (1.0, 1.0);
   (RCLK *> RDATA[13]) = (1.0, 1.0);
   (RCLK *> RDATA[14]) = (1.0, 1.0);
   (RCLK *> RDATA[15]) = (1.0, 1.0);
   $setup(posedge MASK[0], posedge WCLKN, 1.0);
   $setup(negedge MASK[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[0], 1.0);
   $hold(posedge WCLKN, negedge MASK[0], 1.0);
   $setup(posedge MASK[1], posedge WCLKN, 1.0);
   $setup(negedge MASK[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[1], 1.0);
   $hold(posedge WCLKN, negedge MASK[1], 1.0);
   $setup(posedge MASK[2], posedge WCLKN, 1.0);
   $setup(negedge MASK[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[2], 1.0);
   $hold(posedge WCLKN, negedge MASK[2], 1.0);
   $setup(posedge MASK[3], posedge WCLKN, 1.0);
   $setup(negedge MASK[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[3], 1.0);
   $hold(posedge WCLKN, negedge MASK[3], 1.0);
   $setup(posedge MASK[4], posedge WCLKN, 1.0);
   $setup(negedge MASK[4], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[4], 1.0);
   $hold(posedge WCLKN, negedge MASK[4], 1.0);
   $setup(posedge MASK[5], posedge WCLKN, 1.0);
   $setup(negedge MASK[5], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[5], 1.0);
   $hold(posedge WCLKN, negedge MASK[5], 1.0);
   $setup(posedge MASK[6], posedge WCLKN, 1.0);
   $setup(negedge MASK[6], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[6], 1.0);
   $hold(posedge WCLKN, negedge MASK[6], 1.0);
   $setup(posedge MASK[7], posedge WCLKN, 1.0);
   $setup(negedge MASK[7], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[7], 1.0);
   $hold(posedge WCLKN, negedge MASK[7], 1.0);
   $setup(posedge MASK[8], posedge WCLKN, 1.0);
   $setup(negedge MASK[8], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[8], 1.0);
   $hold(posedge WCLKN, negedge MASK[8], 1.0);
   $setup(posedge MASK[9], posedge WCLKN, 1.0);
   $setup(negedge MASK[9], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[9], 1.0);
   $hold(posedge WCLKN, negedge MASK[9], 1.0);
   $setup(posedge MASK[10], posedge WCLKN, 1.0);
   $setup(negedge MASK[10], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[10], 1.0);
   $hold(posedge WCLKN, negedge MASK[10], 1.0);
   $setup(posedge MASK[11], posedge WCLKN, 1.0);
   $setup(negedge MASK[11], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[11], 1.0);
   $hold(posedge WCLKN, negedge MASK[11], 1.0);
   $setup(posedge MASK[12], posedge WCLKN, 1.0);
   $setup(negedge MASK[12], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[12], 1.0);
   $hold(posedge WCLKN, negedge MASK[12], 1.0);
   $setup(posedge MASK[13], posedge WCLKN, 1.0);
   $setup(negedge MASK[13], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[13], 1.0);
   $hold(posedge WCLKN, negedge MASK[13], 1.0);
   $setup(posedge MASK[14], posedge WCLKN, 1.0);
   $setup(negedge MASK[14], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[14], 1.0);
   $hold(posedge WCLKN, negedge MASK[14], 1.0);
   $setup(posedge MASK[15], posedge WCLKN, 1.0);
   $setup(negedge MASK[15], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[15], 1.0);
   $hold(posedge WCLKN, negedge MASK[15], 1.0);
   $setup(posedge WADDR[0], posedge WCLKN, 1.0);
   $setup(negedge WADDR[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[0], 1.0);
   $hold(posedge WCLKN, negedge WADDR[0], 1.0);
   $setup(posedge WADDR[1], posedge WCLKN, 1.0);
   $setup(negedge WADDR[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[1], 1.0);
   $hold(posedge WCLKN, negedge WADDR[1], 1.0);
   $setup(posedge WADDR[2], posedge WCLKN, 1.0);
   $setup(negedge WADDR[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[2], 1.0);
   $hold(posedge WCLKN, negedge WADDR[2], 1.0);
   $setup(posedge WADDR[3], posedge WCLKN, 1.0);
   $setup(negedge WADDR[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[3], 1.0);
   $hold(posedge WCLKN, negedge WADDR[3], 1.0);
   $setup(posedge WADDR[4], posedge WCLKN, 1.0);
   $setup(negedge WADDR[4], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[4], 1.0);
   $hold(posedge WCLKN, negedge WADDR[4], 1.0);
   $setup(posedge WADDR[5], posedge WCLKN, 1.0);
   $setup(negedge WADDR[5], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[5], 1.0);
   $hold(posedge WCLKN, negedge WADDR[5], 1.0);
   $setup(posedge WADDR[6], posedge WCLKN, 1.0);
   $setup(negedge WADDR[6], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[6], 1.0);
   $hold(posedge WCLKN, negedge WADDR[6], 1.0);
   $setup(posedge WADDR[7], posedge WCLKN, 1.0);
   $setup(negedge WADDR[7], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[7], 1.0);
   $hold(posedge WCLKN, negedge WADDR[7], 1.0);
   $setup(posedge WADDR[8], posedge WCLKN, 1.0);
   $setup(negedge WADDR[8], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[8], 1.0);
   $hold(posedge WCLKN, negedge WADDR[8], 1.0);
   $setup(posedge WADDR[9], posedge WCLKN, 1.0);
   $setup(negedge WADDR[9], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[9], 1.0);
   $hold(posedge WCLKN, negedge WADDR[9], 1.0);
   $setup(posedge WDATA[0], posedge WCLKN, 1.0);
   $setup(negedge WDATA[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[0], 1.0);
   $hold(posedge WCLKN, negedge WDATA[0], 1.0);
   $setup(posedge WDATA[1], posedge WCLKN, 1.0);
   $setup(negedge WDATA[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[1], 1.0);
   $hold(posedge WCLKN, negedge WDATA[1], 1.0);
   $setup(posedge WDATA[2], posedge WCLKN, 1.0);
   $setup(negedge WDATA[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[2], 1.0);
   $hold(posedge WCLKN, negedge WDATA[2], 1.0);
   $setup(posedge WDATA[3], posedge WCLKN, 1.0);
   $setup(negedge WDATA[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[3], 1.0);
   $hold(posedge WCLKN, negedge WDATA[3], 1.0);
   $setup(posedge WDATA[4], posedge WCLKN, 1.0);
   $setup(negedge WDATA[4], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[4], 1.0);
   $hold(posedge WCLKN, negedge WDATA[4], 1.0);
   $setup(posedge WDATA[5], posedge WCLKN, 1.0);
   $setup(negedge WDATA[5], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[5], 1.0);
   $hold(posedge WCLKN, negedge WDATA[5], 1.0);
   $setup(posedge WDATA[6], posedge WCLKN, 1.0);
   $setup(negedge WDATA[6], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[6], 1.0);
   $hold(posedge WCLKN, negedge WDATA[6], 1.0);
   $setup(posedge WDATA[7], posedge WCLKN, 1.0);
   $setup(negedge WDATA[7], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[7], 1.0);
   $hold(posedge WCLKN, negedge WDATA[7], 1.0);
   $setup(posedge WDATA[8], posedge WCLKN, 1.0);
   $setup(negedge WDATA[8], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[8], 1.0);
   $hold(posedge WCLKN, negedge WDATA[8], 1.0);
   $setup(posedge WDATA[9], posedge WCLKN, 1.0);
   $setup(negedge WDATA[9], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[9], 1.0);
   $hold(posedge WCLKN, negedge WDATA[9], 1.0);
   $setup(posedge WDATA[10], posedge WCLKN, 1.0);
   $setup(negedge WDATA[10], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[10], 1.0);
   $hold(posedge WCLKN, negedge WDATA[10], 1.0);
   $setup(posedge WDATA[11], posedge WCLKN, 1.0);
   $setup(negedge WDATA[11], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[11], 1.0);
   $hold(posedge WCLKN, negedge WDATA[11], 1.0);
   $setup(posedge WDATA[12], posedge WCLKN, 1.0);
   $setup(negedge WDATA[12], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[12], 1.0);
   $hold(posedge WCLKN, negedge WDATA[12], 1.0);
   $setup(posedge WDATA[13], posedge WCLKN, 1.0);
   $setup(negedge WDATA[13], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[13], 1.0);
   $hold(posedge WCLKN, negedge WDATA[13], 1.0);
   $setup(posedge WDATA[14], posedge WCLKN, 1.0);
   $setup(negedge WDATA[14], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[14], 1.0);
   $hold(posedge WCLKN, negedge WDATA[14], 1.0);
   $setup(posedge WDATA[15], posedge WCLKN, 1.0);
   $setup(negedge WDATA[15], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[15], 1.0);
   $hold(posedge WCLKN, negedge WDATA[15], 1.0);
   $setup(posedge WCLKE, posedge WCLKN, 1.0);
   $setup(negedge WCLKE, posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WCLKE, 1.0);
   $hold(posedge WCLKN, negedge WCLKE, 1.0);
   $setup(posedge WE, posedge WCLKN, 1.0);
   $setup(negedge WE, posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WE, 1.0);
   $hold(posedge WCLKN, negedge WE, 1.0);
   $setup(posedge RADDR[0], posedge RCLK, 1.0);
   $setup(negedge RADDR[0], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[0], 1.0);
   $hold(posedge RCLK, negedge RADDR[0], 1.0);
   $setup(posedge RADDR[1], posedge RCLK, 1.0);
   $setup(negedge RADDR[1], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[1], 1.0);
   $hold(posedge RCLK, negedge RADDR[1], 1.0);
   $setup(posedge RADDR[2], posedge RCLK, 1.0);
   $setup(negedge RADDR[2], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[2], 1.0);
   $hold(posedge RCLK, negedge RADDR[2], 1.0);
   $setup(posedge RADDR[3], posedge RCLK, 1.0);
   $setup(negedge RADDR[3], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[3], 1.0);
   $hold(posedge RCLK, negedge RADDR[3], 1.0);
   $setup(posedge RADDR[4], posedge RCLK, 1.0);
   $setup(negedge RADDR[4], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[4], 1.0);
   $hold(posedge RCLK, negedge RADDR[4], 1.0);
   $setup(posedge RADDR[5], posedge RCLK, 1.0);
   $setup(negedge RADDR[5], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[5], 1.0);
   $hold(posedge RCLK, negedge RADDR[5], 1.0);
   $setup(posedge RADDR[6], posedge RCLK, 1.0);
   $setup(negedge RADDR[6], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[6], 1.0);
   $hold(posedge RCLK, negedge RADDR[6], 1.0);
   $setup(posedge RADDR[7], posedge RCLK, 1.0);
   $setup(negedge RADDR[7], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[7], 1.0);
   $hold(posedge RCLK, negedge RADDR[7], 1.0);
   $setup(posedge RADDR[8], posedge RCLK, 1.0);
   $setup(negedge RADDR[8], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[8], 1.0);
   $hold(posedge RCLK, negedge RADDR[8], 1.0);
   $setup(posedge RADDR[9], posedge RCLK, 1.0);
   $setup(negedge RADDR[9], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[9], 1.0);
   $hold(posedge RCLK, negedge RADDR[9], 1.0);
   $setup(posedge RCLKE, posedge RCLK, 1.0);
   $setup(negedge RCLKE, posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RCLKE, 1.0);
   $hold(posedge RCLK, negedge RCLKE, 1.0);
   $setup(posedge RE, posedge RCLK, 1.0);
   $setup(negedge RE, posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RE, 1.0);
   $hold(posedge RCLK, negedge RE, 1.0);
endspecify
`endif
 
endmodule  // SB_RAM1024x16NW 

//---------------------------------------
//	--- SB_RAM1024x16NRNW -- 
//---------------------------------------
`timescale 1ps/1ps
module SB_RAM1024x16NRNW  ( RDATA, RCLKN, RCLKE, RE, RADDR, WCLKN, WCLKE, WE, WADDR, MASK, WDATA );  

output	[15:0]	RDATA;  
input         	RCLKN;   
input           RCLKE; 
input           RE; 
input	[9:0]   RADDR; 
input           WCLKN; 
input           WCLKE; 
input           WE; 
input 	[9:0]   WADDR; 
input	[15:0]	MASK; 
input 	[15:0]	WDATA; 

parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

wire RCLK, WCLK;
assign (weak0, weak1) RCLKE =1'b1 ;
assign (weak0, weak1) RE =1'b0 ;
assign (weak0, weak1) WCLKE =1'b1 ;
assign (weak0, weak1) WE =1'b0 ;
assign RCLK = ~RCLKN;
assign WCLK = ~WCLKN;

SB_RAM1024x16 sb_ram1024x16rw_inst (
	.RDATA(RDATA),
	.RCLK(RCLK),
	.RCLKE(RCLKE),
	.RE(RE),
	.RADDR(RADDR),
	.WCLK(WCLK),
	.WCLKE(WCLKE),
	.WE(WE),
	.WADDR(WADDR),
	.MASK(MASK),
	.WDATA(WDATA));

defparam sb_ram1024x16rw_inst.INIT_0 = INIT_0;
defparam sb_ram1024x16rw_inst.INIT_1 = INIT_1;
defparam sb_ram1024x16rw_inst.INIT_2 = INIT_2;
defparam sb_ram1024x16rw_inst.INIT_3 = INIT_3;
defparam sb_ram1024x16rw_inst.INIT_4 = INIT_4;
defparam sb_ram1024x16rw_inst.INIT_5 = INIT_5;
defparam sb_ram1024x16rw_inst.INIT_6 = INIT_6;
defparam sb_ram1024x16rw_inst.INIT_7 = INIT_7;
defparam sb_ram1024x16rw_inst.INIT_8 = INIT_8;
defparam sb_ram1024x16rw_inst.INIT_9 = INIT_9;
defparam sb_ram1024x16rw_inst.INIT_A = INIT_A;
defparam sb_ram1024x16rw_inst.INIT_B = INIT_B;
defparam sb_ram1024x16rw_inst.INIT_C = INIT_C;
defparam sb_ram1024x16rw_inst.INIT_D = INIT_D;
defparam sb_ram1024x16rw_inst.INIT_E = INIT_E;
defparam sb_ram1024x16rw_inst.INIT_F = INIT_F;

defparam sb_ram1024x16rw_inst.INIT_10 = INIT_10;
defparam sb_ram1024x16rw_inst.INIT_11 = INIT_11;
defparam sb_ram1024x16rw_inst.INIT_12 = INIT_12;
defparam sb_ram1024x16rw_inst.INIT_13 = INIT_13;
defparam sb_ram1024x16rw_inst.INIT_14 = INIT_14;
defparam sb_ram1024x16rw_inst.INIT_15 = INIT_15;
defparam sb_ram1024x16rw_inst.INIT_16 = INIT_16;
defparam sb_ram1024x16rw_inst.INIT_17 = INIT_17;
defparam sb_ram1024x16rw_inst.INIT_18 = INIT_18;
defparam sb_ram1024x16rw_inst.INIT_19 = INIT_19;
defparam sb_ram1024x16rw_inst.INIT_1A = INIT_1A;
defparam sb_ram1024x16rw_inst.INIT_1B = INIT_1B;
defparam sb_ram1024x16rw_inst.INIT_1C = INIT_1C;
defparam sb_ram1024x16rw_inst.INIT_1D = INIT_1D;
defparam sb_ram1024x16rw_inst.INIT_1E = INIT_1E;
defparam sb_ram1024x16rw_inst.INIT_1F = INIT_1F;

defparam sb_ram1024x16rw_inst.INIT_20 = INIT_20;
defparam sb_ram1024x16rw_inst.INIT_21 = INIT_21;
defparam sb_ram1024x16rw_inst.INIT_22 = INIT_22;
defparam sb_ram1024x16rw_inst.INIT_23 = INIT_23;
defparam sb_ram1024x16rw_inst.INIT_24 = INIT_24;
defparam sb_ram1024x16rw_inst.INIT_25 = INIT_25;
defparam sb_ram1024x16rw_inst.INIT_26 = INIT_26;
defparam sb_ram1024x16rw_inst.INIT_27 = INIT_27;
defparam sb_ram1024x16rw_inst.INIT_28 = INIT_28;
defparam sb_ram1024x16rw_inst.INIT_29 = INIT_29;
defparam sb_ram1024x16rw_inst.INIT_2A = INIT_2A;
defparam sb_ram1024x16rw_inst.INIT_2B = INIT_2B;
defparam sb_ram1024x16rw_inst.INIT_2C = INIT_2C;
defparam sb_ram1024x16rw_inst.INIT_2D = INIT_2D;
defparam sb_ram1024x16rw_inst.INIT_2E = INIT_2E;
defparam sb_ram1024x16rw_inst.INIT_2F = INIT_2F;

defparam sb_ram1024x16rw_inst.INIT_30 = INIT_30;
defparam sb_ram1024x16rw_inst.INIT_31 = INIT_31;
defparam sb_ram1024x16rw_inst.INIT_32 = INIT_32;
defparam sb_ram1024x16rw_inst.INIT_33 = INIT_33;
defparam sb_ram1024x16rw_inst.INIT_34 = INIT_34;
defparam sb_ram1024x16rw_inst.INIT_35 = INIT_35;
defparam sb_ram1024x16rw_inst.INIT_36 = INIT_36;
defparam sb_ram1024x16rw_inst.INIT_37 = INIT_37;
defparam sb_ram1024x16rw_inst.INIT_38 = INIT_38;
defparam sb_ram1024x16rw_inst.INIT_39 = INIT_39;
defparam sb_ram1024x16rw_inst.INIT_3A = INIT_3A;
defparam sb_ram1024x16rw_inst.INIT_3B = INIT_3B;
defparam sb_ram1024x16rw_inst.INIT_3C = INIT_3C;
defparam sb_ram1024x16rw_inst.INIT_3D = INIT_3D;
defparam sb_ram1024x16rw_inst.INIT_3E = INIT_3E;
defparam sb_ram1024x16rw_inst.INIT_3F = INIT_3F;

`ifdef TIMINGCHECK
specify
   (RCLKN *> RDATA[0]) = (1.0, 1.0);
   (RCLKN *> RDATA[1]) = (1.0, 1.0);
   (RCLKN *> RDATA[2]) = (1.0, 1.0);
   (RCLKN *> RDATA[3]) = (1.0, 1.0);
   (RCLKN *> RDATA[4]) = (1.0, 1.0);
   (RCLKN *> RDATA[5]) = (1.0, 1.0);
   (RCLKN *> RDATA[6]) = (1.0, 1.0);
   (RCLKN *> RDATA[7]) = (1.0, 1.0);
   (RCLKN *> RDATA[8]) = (1.0, 1.0);
   (RCLKN *> RDATA[9]) = (1.0, 1.0);
   (RCLKN *> RDATA[10]) = (1.0, 1.0);
   (RCLKN *> RDATA[11]) = (1.0, 1.0);
   (RCLKN *> RDATA[12]) = (1.0, 1.0);
   (RCLKN *> RDATA[13]) = (1.0, 1.0);
   (RCLKN *> RDATA[14]) = (1.0, 1.0);
   (RCLKN *> RDATA[15]) = (1.0, 1.0);
   $setup(posedge MASK[0], posedge WCLKN, 1.0);
   $setup(negedge MASK[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[0], 1.0);
   $hold(posedge WCLKN, negedge MASK[0], 1.0);
   $setup(posedge MASK[1], posedge WCLKN, 1.0);
   $setup(negedge MASK[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[1], 1.0);
   $hold(posedge WCLKN, negedge MASK[1], 1.0);
   $setup(posedge MASK[2], posedge WCLKN, 1.0);
   $setup(negedge MASK[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[2], 1.0);
   $hold(posedge WCLKN, negedge MASK[2], 1.0);
   $setup(posedge MASK[3], posedge WCLKN, 1.0);
   $setup(negedge MASK[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[3], 1.0);
   $hold(posedge WCLKN, negedge MASK[3], 1.0);
   $setup(posedge MASK[4], posedge WCLKN, 1.0);
   $setup(negedge MASK[4], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[4], 1.0);
   $hold(posedge WCLKN, negedge MASK[4], 1.0);
   $setup(posedge MASK[5], posedge WCLKN, 1.0);
   $setup(negedge MASK[5], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[5], 1.0);
   $hold(posedge WCLKN, negedge MASK[5], 1.0);
   $setup(posedge MASK[6], posedge WCLKN, 1.0);
   $setup(negedge MASK[6], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[6], 1.0);
   $hold(posedge WCLKN, negedge MASK[6], 1.0);
   $setup(posedge MASK[7], posedge WCLKN, 1.0);
   $setup(negedge MASK[7], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[7], 1.0);
   $hold(posedge WCLKN, negedge MASK[7], 1.0);
   $setup(posedge MASK[8], posedge WCLKN, 1.0);
   $setup(negedge MASK[8], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[8], 1.0);
   $hold(posedge WCLKN, negedge MASK[8], 1.0);
   $setup(posedge MASK[9], posedge WCLKN, 1.0);
   $setup(negedge MASK[9], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[9], 1.0);
   $hold(posedge WCLKN, negedge MASK[9], 1.0);
   $setup(posedge MASK[10], posedge WCLKN, 1.0);
   $setup(negedge MASK[10], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[10], 1.0);
   $hold(posedge WCLKN, negedge MASK[10], 1.0);
   $setup(posedge MASK[11], posedge WCLKN, 1.0);
   $setup(negedge MASK[11], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[11], 1.0);
   $hold(posedge WCLKN, negedge MASK[11], 1.0);
   $setup(posedge MASK[12], posedge WCLKN, 1.0);
   $setup(negedge MASK[12], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[12], 1.0);
   $hold(posedge WCLKN, negedge MASK[12], 1.0);
   $setup(posedge MASK[13], posedge WCLKN, 1.0);
   $setup(negedge MASK[13], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[13], 1.0);
   $hold(posedge WCLKN, negedge MASK[13], 1.0);
   $setup(posedge MASK[14], posedge WCLKN, 1.0);
   $setup(negedge MASK[14], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[14], 1.0);
   $hold(posedge WCLKN, negedge MASK[14], 1.0);
   $setup(posedge MASK[15], posedge WCLKN, 1.0);
   $setup(negedge MASK[15], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[15], 1.0);
   $hold(posedge WCLKN, negedge MASK[15], 1.0);
   $setup(posedge WADDR[0], posedge WCLKN, 1.0);
   $setup(negedge WADDR[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[0], 1.0);
   $hold(posedge WCLKN, negedge WADDR[0], 1.0);
   $setup(posedge WADDR[1], posedge WCLKN, 1.0);
   $setup(negedge WADDR[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[1], 1.0);
   $hold(posedge WCLKN, negedge WADDR[1], 1.0);
   $setup(posedge WADDR[2], posedge WCLKN, 1.0);
   $setup(negedge WADDR[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[2], 1.0);
   $hold(posedge WCLKN, negedge WADDR[2], 1.0);
   $setup(posedge WADDR[3], posedge WCLKN, 1.0);
   $setup(negedge WADDR[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[3], 1.0);
   $hold(posedge WCLKN, negedge WADDR[3], 1.0);
   $setup(posedge WADDR[4], posedge WCLKN, 1.0);
   $setup(negedge WADDR[4], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[4], 1.0);
   $hold(posedge WCLKN, negedge WADDR[4], 1.0);
   $setup(posedge WADDR[5], posedge WCLKN, 1.0);
   $setup(negedge WADDR[5], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[5], 1.0);
   $hold(posedge WCLKN, negedge WADDR[5], 1.0);
   $setup(posedge WADDR[6], posedge WCLKN, 1.0);
   $setup(negedge WADDR[6], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[6], 1.0);
   $hold(posedge WCLKN, negedge WADDR[6], 1.0);
   $setup(posedge WADDR[7], posedge WCLKN, 1.0);
   $setup(negedge WADDR[7], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[7], 1.0);
   $hold(posedge WCLKN, negedge WADDR[7], 1.0);
   $setup(posedge WADDR[8], posedge WCLKN, 1.0);
   $setup(negedge WADDR[8], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[8], 1.0);
   $hold(posedge WCLKN, negedge WADDR[8], 1.0);
   $setup(posedge WADDR[9], posedge WCLKN, 1.0);
   $setup(negedge WADDR[9], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[9], 1.0);
   $hold(posedge WCLKN, negedge WADDR[9], 1.0);
   $setup(posedge WDATA[0], posedge WCLKN, 1.0);
   $setup(negedge WDATA[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[0], 1.0);
   $hold(posedge WCLKN, negedge WDATA[0], 1.0);
   $setup(posedge WDATA[1], posedge WCLKN, 1.0);
   $setup(negedge WDATA[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[1], 1.0);
   $hold(posedge WCLKN, negedge WDATA[1], 1.0);
   $setup(posedge WDATA[2], posedge WCLKN, 1.0);
   $setup(negedge WDATA[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[2], 1.0);
   $hold(posedge WCLKN, negedge WDATA[2], 1.0);
   $setup(posedge WDATA[3], posedge WCLKN, 1.0);
   $setup(negedge WDATA[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[3], 1.0);
   $hold(posedge WCLKN, negedge WDATA[3], 1.0);
   $setup(posedge WDATA[4], posedge WCLKN, 1.0);
   $setup(negedge WDATA[4], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[4], 1.0);
   $hold(posedge WCLKN, negedge WDATA[4], 1.0);
   $setup(posedge WDATA[5], posedge WCLKN, 1.0);
   $setup(negedge WDATA[5], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[5], 1.0);
   $hold(posedge WCLKN, negedge WDATA[5], 1.0);
   $setup(posedge WDATA[6], posedge WCLKN, 1.0);
   $setup(negedge WDATA[6], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[6], 1.0);
   $hold(posedge WCLKN, negedge WDATA[6], 1.0);
   $setup(posedge WDATA[7], posedge WCLKN, 1.0);
   $setup(negedge WDATA[7], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[7], 1.0);
   $hold(posedge WCLKN, negedge WDATA[7], 1.0);
   $setup(posedge WDATA[8], posedge WCLKN, 1.0);
   $setup(negedge WDATA[8], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[8], 1.0);
   $hold(posedge WCLKN, negedge WDATA[8], 1.0);
   $setup(posedge WDATA[9], posedge WCLKN, 1.0);
   $setup(negedge WDATA[9], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[9], 1.0);
   $hold(posedge WCLKN, negedge WDATA[9], 1.0);
   $setup(posedge WDATA[10], posedge WCLKN, 1.0);
   $setup(negedge WDATA[10], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[10], 1.0);
   $hold(posedge WCLKN, negedge WDATA[10], 1.0);
   $setup(posedge WDATA[11], posedge WCLKN, 1.0);
   $setup(negedge WDATA[11], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[11], 1.0);
   $hold(posedge WCLKN, negedge WDATA[11], 1.0);
   $setup(posedge WDATA[12], posedge WCLKN, 1.0);
   $setup(negedge WDATA[12], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[12], 1.0);
   $hold(posedge WCLKN, negedge WDATA[12], 1.0);
   $setup(posedge WDATA[13], posedge WCLKN, 1.0);
   $setup(negedge WDATA[13], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[13], 1.0);
   $hold(posedge WCLKN, negedge WDATA[13], 1.0);
   $setup(posedge WDATA[14], posedge WCLKN, 1.0);
   $setup(negedge WDATA[14], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[14], 1.0);
   $hold(posedge WCLKN, negedge WDATA[14], 1.0);
   $setup(posedge WDATA[15], posedge WCLKN, 1.0);
   $setup(negedge WDATA[15], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[15], 1.0);
   $hold(posedge WCLKN, negedge WDATA[15], 1.0);
   $setup(posedge WCLKE, posedge WCLKN, 1.0);
   $setup(negedge WCLKE, posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WCLKE, 1.0);
   $hold(posedge WCLKN, negedge WCLKE, 1.0);
   $setup(posedge WE, posedge WCLKN, 1.0);
   $setup(negedge WE, posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WE, 1.0);
   $hold(posedge WCLKN, negedge WE, 1.0);
   $setup(posedge RADDR[0], posedge RCLKN, 1.0);
   $setup(negedge RADDR[0], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[0], 1.0);
   $hold(posedge RCLKN, negedge RADDR[0], 1.0);
   $setup(posedge RADDR[1], posedge RCLKN, 1.0);
   $setup(negedge RADDR[1], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[1], 1.0);
   $hold(posedge RCLKN, negedge RADDR[1], 1.0);
   $setup(posedge RADDR[2], posedge RCLKN, 1.0);
   $setup(negedge RADDR[2], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[2], 1.0);
   $hold(posedge RCLKN, negedge RADDR[2], 1.0);
   $setup(posedge RADDR[3], posedge RCLKN, 1.0);
   $setup(negedge RADDR[3], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[3], 1.0);
   $hold(posedge RCLKN, negedge RADDR[3], 1.0);
   $setup(posedge RADDR[4], posedge RCLKN, 1.0);
   $setup(negedge RADDR[4], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[4], 1.0);
   $hold(posedge RCLKN, negedge RADDR[4], 1.0);
   $setup(posedge RADDR[5], posedge RCLKN, 1.0);
   $setup(negedge RADDR[5], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[5], 1.0);
   $hold(posedge RCLKN, negedge RADDR[5], 1.0);
   $setup(posedge RADDR[6], posedge RCLKN, 1.0);
   $setup(negedge RADDR[6], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[6], 1.0);
   $hold(posedge RCLKN, negedge RADDR[6], 1.0);
   $setup(posedge RADDR[7], posedge RCLKN, 1.0);
   $setup(negedge RADDR[7], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[7], 1.0);
   $hold(posedge RCLKN, negedge RADDR[7], 1.0);
   $setup(posedge RADDR[8], posedge RCLKN, 1.0);
   $setup(negedge RADDR[8], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[8], 1.0);
   $hold(posedge RCLKN, negedge RADDR[8], 1.0);
   $setup(posedge RADDR[9], posedge RCLKN, 1.0);
   $setup(negedge RADDR[9], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[9], 1.0);
   $hold(posedge RCLKN, negedge RADDR[9], 1.0);
   $setup(posedge RCLKE, posedge RCLKN, 1.0);
   $setup(negedge RCLKE, posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RCLKE, 1.0);
   $hold(posedge RCLKN, negedge RCLKE, 1.0);
   $setup(posedge RE, posedge RCLKN, 1.0);
   $setup(negedge RE, posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RE, 1.0);
   $hold(posedge RCLKN, negedge RE, 1.0);
endspecify
`endif

endmodule  // SB_RAM1024x16NRNW

//---------------------------------------
//	--- SB_RAM2048x8
//---------------------------------------
`timescale 1ps/1ps
module SB_RAM2048x8 (RDATA, RCLK, RCLKE, RE, RADDR, WCLK, WCLKE, WE, WADDR, WDATA ); 

output	[7:0]	RDATA;  
input         	RCLK;   
input           RCLKE; 
input           RE; 
input	[10:0]  RADDR; 
input           WCLK; 
input           WCLKE; 
input           WE; 
input 	[10:0]  WADDR; 
input 	[7:0]	WDATA; 

parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;


// local Parameters
localparam			CLOCK_PERIOD = 200;	//
localparam 			DELAY	= (CLOCK_PERIOD/10);		// Clock-to-output delay. Zero
							// time delays can be confusing
							// and sometimes cause problems.
localparam 			BUS_WIDTH = 8;		// Width of RAM (number of bits)

localparam 			ADDRESS_BUS_SIZE = 11;	// Number of bits required to
							// represent the RAM address

localparam   ADDRESSABLE_SPACE  = 2**ADDRESS_BUS_SIZE;	// Decimal address range [2^Size:0]


// SIGNAL DECLARATIONS
wire			   	WCLK_g, RCLK_g;
reg 				WCLKE_sync, RCLKE_sync; 
assign (weak0, weak1) RCLKE =1'b1 ;
assign (weak0, weak1) RE =1'b0 ;
assign (weak0, weak1) WCLKE =1'b1 ;
assign (weak0, weak1) WE =1'b0 ;
reg	Memory	[BUS_WIDTH*ADDRESSABLE_SPACE-1:0];
// 
event Read_e, Write_e;

//////////////////// Collision detect begins here ///////////////////////////////
localparam 	TRUE = 1'b1;
localparam	FALSE = 1'b0;
reg 		Time_Collision_Detected = 1'b0;
wire		Address_Collision_Detected;

event Collision_e;

time COLLISION_TIME_WINDOW = (CLOCK_PERIOD/8); // This is an arbitray value, but is better than using an absolute 
						    // value, because the actual time window depends on the actual silicon 
						    // implementation. Thus the test is indicative of an Error and not
						    // guaranteed to be an error. Even so this is usefull.
time time_WCLK_RCLK, time_WCLK, time_RCLK;


//function reg Check_Timed_Window_Violation;
function	Check_Timed_Window_Violation;	
input T1, T2, Minimum_Time_Window;
time T1, T2;
time Minimum_Time_Window;
time Difference;	
	begin
		Difference = (T1 - T2);
		if (Difference < 0) Difference = -Difference;
		Check_Timed_Window_Violation = (Difference < Minimum_Time_Window);
	end
endfunction


initial begin
       time_WCLK = CLOCK_PERIOD;	// Arbitrary initialisation value, ensure no window collison error on first clock edge.
       time_RCLK = (CLOCK_PERIOD*8);	// Arbitrary initialisation difference value, ensure no collision error on first clock edge.					
end

integer	i,j;


initial	//	initialize ram_16k (2048 x 8) by init  parameters, section by section
begin
	for	(i=0; i<=(256/BUS_WIDTH)-1; i=i+1)       
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)    
		begin 
			Memory[BUS_WIDTH*i+j]		=	INIT_0[BUS_WIDTH*i+j];
			Memory[256*1+BUS_WIDTH*i+j]	=	INIT_1[BUS_WIDTH*i+j];
			Memory[256*2+BUS_WIDTH*i+j]	=	INIT_2[BUS_WIDTH*i+j];
			Memory[256*3+BUS_WIDTH*i+j]	=	INIT_3[BUS_WIDTH*i+j];
			Memory[256*4+BUS_WIDTH*i+j]	=	INIT_4[BUS_WIDTH*i+j];
			Memory[256*5+BUS_WIDTH*i+j]	=	INIT_5[BUS_WIDTH*i+j];
			Memory[256*6+BUS_WIDTH*i+j]	=	INIT_6[BUS_WIDTH*i+j];
			Memory[256*7+BUS_WIDTH*i+j]	=	INIT_7[BUS_WIDTH*i+j];
			Memory[256*8+BUS_WIDTH*i+j]	=	INIT_8[BUS_WIDTH*i+j];
			Memory[256*9+BUS_WIDTH*i+j]	=	INIT_9[BUS_WIDTH*i+j];
			Memory[256*10+BUS_WIDTH*i+j]	=	INIT_A[BUS_WIDTH*i+j];
			Memory[256*11+BUS_WIDTH*i+j]	=	INIT_B[BUS_WIDTH*i+j];
			Memory[256*12+BUS_WIDTH*i+j]	=	INIT_C[BUS_WIDTH*i+j];
			Memory[256*13+BUS_WIDTH*i+j]	=	INIT_D[BUS_WIDTH*i+j];
			Memory[256*14+BUS_WIDTH*i+j]	=	INIT_E[BUS_WIDTH*i+j];
			Memory[256*15+BUS_WIDTH*i+j]	=	INIT_F[BUS_WIDTH*i+j];

			Memory[256*16+BUS_WIDTH*i+j]	=	INIT_10[BUS_WIDTH*i+j];
			Memory[256*17+BUS_WIDTH*i+j]	=	INIT_11[BUS_WIDTH*i+j];
			Memory[256*18+BUS_WIDTH*i+j]	=	INIT_12[BUS_WIDTH*i+j];
			Memory[256*19+BUS_WIDTH*i+j]	=	INIT_13[BUS_WIDTH*i+j];
			Memory[256*20+BUS_WIDTH*i+j]	=	INIT_14[BUS_WIDTH*i+j];
			Memory[256*21+BUS_WIDTH*i+j]	=	INIT_15[BUS_WIDTH*i+j];
			Memory[256*22+BUS_WIDTH*i+j]	=	INIT_16[BUS_WIDTH*i+j];
			Memory[256*23+BUS_WIDTH*i+j]	=	INIT_17[BUS_WIDTH*i+j];
			Memory[256*24+BUS_WIDTH*i+j]	=	INIT_18[BUS_WIDTH*i+j];
			Memory[256*25+BUS_WIDTH*i+j]	=	INIT_19[BUS_WIDTH*i+j];
			Memory[256*26+BUS_WIDTH*i+j]	=	INIT_1A[BUS_WIDTH*i+j];
			Memory[256*27+BUS_WIDTH*i+j]	=	INIT_1B[BUS_WIDTH*i+j];
			Memory[256*28+BUS_WIDTH*i+j]	=	INIT_1C[BUS_WIDTH*i+j];
			Memory[256*29+BUS_WIDTH*i+j]	=	INIT_1D[BUS_WIDTH*i+j];
			Memory[256*30+BUS_WIDTH*i+j]	=	INIT_1E[BUS_WIDTH*i+j];
			Memory[256*31+BUS_WIDTH*i+j]	=	INIT_1F[BUS_WIDTH*i+j];

			Memory[256*32+BUS_WIDTH*i+j]	=	INIT_20[BUS_WIDTH*i+j];
			Memory[256*33+BUS_WIDTH*i+j]	=	INIT_21[BUS_WIDTH*i+j];
			Memory[256*34+BUS_WIDTH*i+j]	=	INIT_22[BUS_WIDTH*i+j];
			Memory[256*35+BUS_WIDTH*i+j]	=	INIT_23[BUS_WIDTH*i+j];
			Memory[256*36+BUS_WIDTH*i+j]	=	INIT_24[BUS_WIDTH*i+j];
			Memory[256*37+BUS_WIDTH*i+j]	=	INIT_25[BUS_WIDTH*i+j];
			Memory[256*38+BUS_WIDTH*i+j]	=	INIT_26[BUS_WIDTH*i+j];
			Memory[256*39+BUS_WIDTH*i+j]	=	INIT_27[BUS_WIDTH*i+j];
			Memory[256*40+BUS_WIDTH*i+j]	=	INIT_28[BUS_WIDTH*i+j];
			Memory[256*41+BUS_WIDTH*i+j]	=	INIT_29[BUS_WIDTH*i+j];
			Memory[256*42+BUS_WIDTH*i+j]	=	INIT_2A[BUS_WIDTH*i+j];
			Memory[256*43+BUS_WIDTH*i+j]	=	INIT_2B[BUS_WIDTH*i+j];
			Memory[256*44+BUS_WIDTH*i+j]	=	INIT_2C[BUS_WIDTH*i+j];
			Memory[256*45+BUS_WIDTH*i+j]	=	INIT_2D[BUS_WIDTH*i+j];
			Memory[256*46+BUS_WIDTH*i+j]	=	INIT_2E[BUS_WIDTH*i+j];
			Memory[256*47+BUS_WIDTH*i+j]	=	INIT_2F[BUS_WIDTH*i+j];

			Memory[256*48+BUS_WIDTH*i+j]	=	INIT_30[BUS_WIDTH*i+j];
			Memory[256*49+BUS_WIDTH*i+j]	=	INIT_31[BUS_WIDTH*i+j];
			Memory[256*50+BUS_WIDTH*i+j]	=	INIT_32[BUS_WIDTH*i+j];
			Memory[256*51+BUS_WIDTH*i+j]	=	INIT_33[BUS_WIDTH*i+j];
			Memory[256*52+BUS_WIDTH*i+j]	=	INIT_34[BUS_WIDTH*i+j];
			Memory[256*53+BUS_WIDTH*i+j]	=	INIT_35[BUS_WIDTH*i+j];
			Memory[256*54+BUS_WIDTH*i+j]	=	INIT_36[BUS_WIDTH*i+j];
			Memory[256*55+BUS_WIDTH*i+j]	=	INIT_37[BUS_WIDTH*i+j];
			Memory[256*56+BUS_WIDTH*i+j]	=	INIT_38[BUS_WIDTH*i+j];
			Memory[256*57+BUS_WIDTH*i+j]	=	INIT_39[BUS_WIDTH*i+j];
			Memory[256*58+BUS_WIDTH*i+j]	=	INIT_3A[BUS_WIDTH*i+j];
			Memory[256*59+BUS_WIDTH*i+j]	=	INIT_3B[BUS_WIDTH*i+j];
			Memory[256*60+BUS_WIDTH*i+j]	=	INIT_3C[BUS_WIDTH*i+j];
			Memory[256*61+BUS_WIDTH*i+j]	=	INIT_3D[BUS_WIDTH*i+j];
			Memory[256*62+BUS_WIDTH*i+j]	=	INIT_3E[BUS_WIDTH*i+j];
			Memory[256*63+BUS_WIDTH*i+j]	=	INIT_3F[BUS_WIDTH*i+j];
		end 
	end

end

assign Address_Collision_Detected = ((RE & WE & WCLKE & RCLKE)&(WADDR == RADDR)); 

always @(WCLK or WCLKE) 
begin 
	if(~WCLK)
	WCLKE_sync = WCLKE;   	
end 

always @(RCLK or RCLKE) 
begin 
	if (~RCLK)
	RCLKE_sync = RCLKE; 	
end 

assign WCLK_g = WCLK & WCLKE_sync;
assign RCLK_g = RCLK & RCLKE_sync;


always @(posedge WCLK_g) begin
	time_WCLK = $time;
end

always @(posedge RCLK_g) begin
    	time_RCLK = $time;
end
integer	SB_RAM2048x8_RDATA_log_file;					//.....................
initial	SB_RAM2048x8_RDATA_log_file=("SB_RAM2048x8_RDATA_log_file.txt");	//.....................
always @(posedge WCLK_g) begin

	Time_Collision_Detected = Check_Timed_Window_Violation(time_WCLK,time_RCLK,COLLISION_TIME_WINDOW);
        if (Time_Collision_Detected & Address_Collision_Detected)begin
        	$display("Warning: Write-Read collision detected, Data read value is XXXX\n");
 		$display("WCLK Time: %.3f   RCLK Time:%.3f  ",time_WCLK, time_RCLK,"WADDR: %d   RADDR:%d\n",WADDR, RADDR); 
 		$fdisplay(SB_RAM2048x8_RDATA_log_file,"Warning: Write-Read collision detected, Data read value is XXXX\n");
		$fdisplay(SB_RAM2048x8_RDATA_log_file,"WCLK Time: %.3f   RCLK Time:%.3f  ",time_WCLK, time_RCLK, "WADDR: %d   RADDR:%d\n",WADDR, RADDR); 	
 		-> Collision_e;
	end
end

//	code modify for universal verilog compiler

always @ (posedge WCLK_g)
begin
	if	(WE)
	begin
		-> Write_e;
		for	(i=0;i<=BUS_WIDTH-1; i=i+1)
		begin
				Memory[WADDR*BUS_WIDTH+i]	<=	WDATA[i];
		end
	end
end

reg	[BUS_WIDTH-1:0]	RDATA = 0;

// Look at the rising edge of the clock

always @ (posedge RCLK_g)
begin
	if	(RE)
	begin
		-> Read_e;
		if	(Time_Collision_Detected & Address_Collision_Detected) 
			RDATA <= {BUS_WIDTH{1'hX}};
		else
			for	(i=0;i<=BUS_WIDTH-1;i=i+1)
				RDATA[i]	<= Memory[RADDR*BUS_WIDTH+i];
	end
end

`ifdef TIMINGCHECK
specify
   (RCLK *> RDATA[0]) = (1.0, 1.0);
   (RCLK *> RDATA[1]) = (1.0, 1.0);
   (RCLK *> RDATA[2]) = (1.0, 1.0);
   (RCLK *> RDATA[3]) = (1.0, 1.0);
   (RCLK *> RDATA[4]) = (1.0, 1.0);
   (RCLK *> RDATA[5]) = (1.0, 1.0);
   (RCLK *> RDATA[6]) = (1.0, 1.0);
   (RCLK *> RDATA[7]) = (1.0, 1.0);
   $setup(posedge WADDR[0], posedge WCLK, 1.0);
   $setup(negedge WADDR[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[0], 1.0);
   $hold(posedge WCLK, negedge WADDR[0], 1.0);
   $setup(posedge WADDR[1], posedge WCLK, 1.0);
   $setup(negedge WADDR[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[1], 1.0);
   $hold(posedge WCLK, negedge WADDR[1], 1.0);
   $setup(posedge WADDR[2], posedge WCLK, 1.0);
   $setup(negedge WADDR[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[2], 1.0);
   $hold(posedge WCLK, negedge WADDR[2], 1.0);
   $setup(posedge WADDR[3], posedge WCLK, 1.0);
   $setup(negedge WADDR[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[3], 1.0);
   $hold(posedge WCLK, negedge WADDR[3], 1.0);
   $setup(posedge WADDR[4], posedge WCLK, 1.0);
   $setup(negedge WADDR[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[4], 1.0);
   $hold(posedge WCLK, negedge WADDR[4], 1.0);
   $setup(posedge WADDR[5], posedge WCLK, 1.0);
   $setup(negedge WADDR[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[5], 1.0);
   $hold(posedge WCLK, negedge WADDR[5], 1.0);
   $setup(posedge WADDR[6], posedge WCLK, 1.0);
   $setup(negedge WADDR[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[6], 1.0);
   $hold(posedge WCLK, negedge WADDR[6], 1.0);
   $setup(posedge WADDR[7], posedge WCLK, 1.0);
   $setup(negedge WADDR[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[7], 1.0);
   $hold(posedge WCLK, negedge WADDR[7], 1.0);
   $setup(posedge WADDR[8], posedge WCLK, 1.0);
   $setup(negedge WADDR[8], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[8], 1.0);
   $hold(posedge WCLK, negedge WADDR[8], 1.0);
   $setup(posedge WADDR[9], posedge WCLK, 1.0);
   $setup(negedge WADDR[9], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[9], 1.0);
   $hold(posedge WCLK, negedge WADDR[9], 1.0);
   $setup(posedge WADDR[10], posedge WCLK, 1.0);
   $setup(negedge WADDR[10], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[10], 1.0);
   $hold(posedge WCLK, negedge WADDR[10], 1.0);
   $setup(posedge WDATA[0], posedge WCLK, 1.0);
   $setup(negedge WDATA[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[0], 1.0);
   $hold(posedge WCLK, negedge WDATA[0], 1.0);
   $setup(posedge WDATA[1], posedge WCLK, 1.0);
   $setup(negedge WDATA[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[1], 1.0);
   $hold(posedge WCLK, negedge WDATA[1], 1.0);
   $setup(posedge WDATA[2], posedge WCLK, 1.0);
   $setup(negedge WDATA[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[2], 1.0);
   $hold(posedge WCLK, negedge WDATA[2], 1.0);
   $setup(posedge WDATA[3], posedge WCLK, 1.0);
   $setup(negedge WDATA[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[3], 1.0);
   $hold(posedge WCLK, negedge WDATA[3], 1.0);
   $setup(posedge WDATA[4], posedge WCLK, 1.0);
   $setup(negedge WDATA[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[4], 1.0);
   $hold(posedge WCLK, negedge WDATA[4], 1.0);
   $setup(posedge WDATA[5], posedge WCLK, 1.0);
   $setup(negedge WDATA[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[5], 1.0);
   $hold(posedge WCLK, negedge WDATA[5], 1.0);
   $setup(posedge WDATA[6], posedge WCLK, 1.0);
   $setup(negedge WDATA[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[6], 1.0);
   $hold(posedge WCLK, negedge WDATA[6], 1.0);
   $setup(posedge WDATA[7], posedge WCLK, 1.0);
   $setup(negedge WDATA[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[7], 1.0);
   $hold(posedge WCLK, negedge WDATA[7], 1.0);
   $setup(posedge WCLKE, posedge WCLK, 1.0);
   $setup(negedge WCLKE, posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WCLKE, 1.0);
   $hold(posedge WCLK, negedge WCLKE, 1.0);
   $setup(posedge WE, posedge WCLK, 1.0);
   $setup(negedge WE, posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WE, 1.0);
   $hold(posedge WCLK, negedge WE, 1.0);
   $setup(posedge RADDR[0], posedge RCLK, 1.0);
   $setup(negedge RADDR[0], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[0], 1.0);
   $hold(posedge RCLK, negedge RADDR[0], 1.0);
   $setup(posedge RADDR[1], posedge RCLK, 1.0);
   $setup(negedge RADDR[1], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[1], 1.0);
   $hold(posedge RCLK, negedge RADDR[1], 1.0);
   $setup(posedge RADDR[2], posedge RCLK, 1.0);
   $setup(negedge RADDR[2], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[2], 1.0);
   $hold(posedge RCLK, negedge RADDR[2], 1.0);
   $setup(posedge RADDR[3], posedge RCLK, 1.0);
   $setup(negedge RADDR[3], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[3], 1.0);
   $hold(posedge RCLK, negedge RADDR[3], 1.0);
   $setup(posedge RADDR[4], posedge RCLK, 1.0);
   $setup(negedge RADDR[4], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[4], 1.0);
   $hold(posedge RCLK, negedge RADDR[4], 1.0);
   $setup(posedge RADDR[5], posedge RCLK, 1.0);
   $setup(negedge RADDR[5], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[5], 1.0);
   $hold(posedge RCLK, negedge RADDR[5], 1.0);
   $setup(posedge RADDR[6], posedge RCLK, 1.0);
   $setup(negedge RADDR[6], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[6], 1.0);
   $hold(posedge RCLK, negedge RADDR[6], 1.0);
   $setup(posedge RADDR[7], posedge RCLK, 1.0);
   $setup(negedge RADDR[7], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[7], 1.0);
   $hold(posedge RCLK, negedge RADDR[7], 1.0);
   $setup(posedge RADDR[8], posedge RCLK, 1.0);
   $setup(negedge RADDR[8], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[8], 1.0);
   $hold(posedge RCLK, negedge RADDR[8], 1.0);
   $setup(posedge RADDR[9], posedge RCLK, 1.0);
   $setup(negedge RADDR[9], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[9], 1.0);
   $hold(posedge RCLK, negedge RADDR[9], 1.0);
   $setup(posedge RADDR[10], posedge RCLK, 1.0);
   $setup(negedge RADDR[10], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[10], 1.0);
   $hold(posedge RCLK, negedge RADDR[10], 1.0);
   $setup(posedge RCLKE, posedge RCLK, 1.0);
   $setup(negedge RCLKE, posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RCLKE, 1.0);
   $hold(posedge RCLK, negedge RCLKE, 1.0);
   $setup(posedge RE, posedge RCLK, 1.0);
   $setup(negedge RE, posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RE, 1.0);
   $hold(posedge RCLK, negedge RE, 1.0);
endspecify
`endif

endmodule //  SB_RAM2048x8

//---------------------------------------
//	--- SB_RAM2048x8NR
//---------------------------------------
`timescale 1ps/1ps
module SB_RAM2048x8NR ( RDATA, RCLKN, RCLKE, RE, RADDR, WCLK, WCLKE, WE, WADDR, WDATA );  

output	[7:0]	RDATA;  
input         	RCLKN;   
input           RCLKE; 
input           RE; 
input	[10:0]  RADDR; 
input           WCLK; 
input           WCLKE; 
input           WE; 
input 	[10:0]  WADDR; 
input 	[7:0]	WDATA; 

parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

wire RCLK;
assign (weak0, weak1) RCLKE =1'b1 ;
assign (weak0, weak1) RE =1'b0 ;
assign (weak0, weak1) WCLKE =1'b1 ;
assign (weak0, weak1) WE =1'b0 ;
assign RCLK = ~RCLKN;

SB_RAM2048x8 sb_ram2048x8r_inst (
	.RDATA(RDATA),
	.RCLK(RCLK),
	.RCLKE(RCLKE),
	.RE(RE),
	.RADDR(RADDR),
	.WCLK(WCLK),
	.WCLKE(WCLKE),
	.WE(WE),
	.WADDR(WADDR),
	.WDATA(WDATA));

defparam sb_ram2048x8r_inst.INIT_0 = INIT_0;
defparam sb_ram2048x8r_inst.INIT_1 = INIT_1;
defparam sb_ram2048x8r_inst.INIT_2 = INIT_2;
defparam sb_ram2048x8r_inst.INIT_3 = INIT_3;
defparam sb_ram2048x8r_inst.INIT_4 = INIT_4;
defparam sb_ram2048x8r_inst.INIT_5 = INIT_5;
defparam sb_ram2048x8r_inst.INIT_6 = INIT_6;
defparam sb_ram2048x8r_inst.INIT_7 = INIT_7;
defparam sb_ram2048x8r_inst.INIT_8 = INIT_8;
defparam sb_ram2048x8r_inst.INIT_9 = INIT_9;
defparam sb_ram2048x8r_inst.INIT_A = INIT_A;
defparam sb_ram2048x8r_inst.INIT_B = INIT_B;
defparam sb_ram2048x8r_inst.INIT_C = INIT_C;
defparam sb_ram2048x8r_inst.INIT_D = INIT_D;
defparam sb_ram2048x8r_inst.INIT_E = INIT_E;
defparam sb_ram2048x8r_inst.INIT_F = INIT_F;

defparam sb_ram2048x8r_inst.INIT_10 = INIT_10;
defparam sb_ram2048x8r_inst.INIT_11 = INIT_11;
defparam sb_ram2048x8r_inst.INIT_12 = INIT_12;
defparam sb_ram2048x8r_inst.INIT_13 = INIT_13;
defparam sb_ram2048x8r_inst.INIT_14 = INIT_14;
defparam sb_ram2048x8r_inst.INIT_15 = INIT_15;
defparam sb_ram2048x8r_inst.INIT_16 = INIT_16;
defparam sb_ram2048x8r_inst.INIT_17 = INIT_17;
defparam sb_ram2048x8r_inst.INIT_18 = INIT_18;
defparam sb_ram2048x8r_inst.INIT_19 = INIT_19;
defparam sb_ram2048x8r_inst.INIT_1A = INIT_1A;
defparam sb_ram2048x8r_inst.INIT_1B = INIT_1B;
defparam sb_ram2048x8r_inst.INIT_1C = INIT_1C;
defparam sb_ram2048x8r_inst.INIT_1D = INIT_1D;
defparam sb_ram2048x8r_inst.INIT_1E = INIT_1E;
defparam sb_ram2048x8r_inst.INIT_1F = INIT_1F;

defparam sb_ram2048x8r_inst.INIT_20 = INIT_20;
defparam sb_ram2048x8r_inst.INIT_21 = INIT_21;
defparam sb_ram2048x8r_inst.INIT_22 = INIT_22;
defparam sb_ram2048x8r_inst.INIT_23 = INIT_23;
defparam sb_ram2048x8r_inst.INIT_24 = INIT_24;
defparam sb_ram2048x8r_inst.INIT_25 = INIT_25;
defparam sb_ram2048x8r_inst.INIT_26 = INIT_26;
defparam sb_ram2048x8r_inst.INIT_27 = INIT_27;
defparam sb_ram2048x8r_inst.INIT_28 = INIT_28;
defparam sb_ram2048x8r_inst.INIT_29 = INIT_29;
defparam sb_ram2048x8r_inst.INIT_2A = INIT_2A;
defparam sb_ram2048x8r_inst.INIT_2B = INIT_2B;
defparam sb_ram2048x8r_inst.INIT_2C = INIT_2C;
defparam sb_ram2048x8r_inst.INIT_2D = INIT_2D;
defparam sb_ram2048x8r_inst.INIT_2E = INIT_2E;
defparam sb_ram2048x8r_inst.INIT_2F = INIT_2F;

defparam sb_ram2048x8r_inst.INIT_30 = INIT_30;
defparam sb_ram2048x8r_inst.INIT_31 = INIT_31;
defparam sb_ram2048x8r_inst.INIT_32 = INIT_32;
defparam sb_ram2048x8r_inst.INIT_33 = INIT_33;
defparam sb_ram2048x8r_inst.INIT_34 = INIT_34;
defparam sb_ram2048x8r_inst.INIT_35 = INIT_35;
defparam sb_ram2048x8r_inst.INIT_36 = INIT_36;
defparam sb_ram2048x8r_inst.INIT_37 = INIT_37;
defparam sb_ram2048x8r_inst.INIT_38 = INIT_38;
defparam sb_ram2048x8r_inst.INIT_39 = INIT_39;
defparam sb_ram2048x8r_inst.INIT_3A = INIT_3A;
defparam sb_ram2048x8r_inst.INIT_3B = INIT_3B;
defparam sb_ram2048x8r_inst.INIT_3C = INIT_3C;
defparam sb_ram2048x8r_inst.INIT_3D = INIT_3D;
defparam sb_ram2048x8r_inst.INIT_3E = INIT_3E;
defparam sb_ram2048x8r_inst.INIT_3F = INIT_3F;


`ifdef TIMINGCHECK
specify
   (RCLKN *> RDATA[0]) = (1.0, 1.0);
   (RCLKN *> RDATA[1]) = (1.0, 1.0);
   (RCLKN *> RDATA[2]) = (1.0, 1.0);
   (RCLKN *> RDATA[3]) = (1.0, 1.0);
   (RCLKN *> RDATA[4]) = (1.0, 1.0);
   (RCLKN *> RDATA[5]) = (1.0, 1.0);
   (RCLKN *> RDATA[6]) = (1.0, 1.0);
   (RCLKN *> RDATA[7]) = (1.0, 1.0);
   $setup(posedge WADDR[0], posedge WCLK, 1.0);
   $setup(negedge WADDR[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[0], 1.0);
   $hold(posedge WCLK, negedge WADDR[0], 1.0);
   $setup(posedge WADDR[1], posedge WCLK, 1.0);
   $setup(negedge WADDR[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[1], 1.0);
   $hold(posedge WCLK, negedge WADDR[1], 1.0);
   $setup(posedge WADDR[2], posedge WCLK, 1.0);
   $setup(negedge WADDR[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[2], 1.0);
   $hold(posedge WCLK, negedge WADDR[2], 1.0);
   $setup(posedge WADDR[3], posedge WCLK, 1.0);
   $setup(negedge WADDR[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[3], 1.0);
   $hold(posedge WCLK, negedge WADDR[3], 1.0);
   $setup(posedge WADDR[4], posedge WCLK, 1.0);
   $setup(negedge WADDR[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[4], 1.0);
   $hold(posedge WCLK, negedge WADDR[4], 1.0);
   $setup(posedge WADDR[5], posedge WCLK, 1.0);
   $setup(negedge WADDR[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[5], 1.0);
   $hold(posedge WCLK, negedge WADDR[5], 1.0);
   $setup(posedge WADDR[6], posedge WCLK, 1.0);
   $setup(negedge WADDR[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[6], 1.0);
   $hold(posedge WCLK, negedge WADDR[6], 1.0);
   $setup(posedge WADDR[7], posedge WCLK, 1.0);
   $setup(negedge WADDR[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[7], 1.0);
   $hold(posedge WCLK, negedge WADDR[7], 1.0);
   $setup(posedge WADDR[8], posedge WCLK, 1.0);
   $setup(negedge WADDR[8], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[8], 1.0);
   $hold(posedge WCLK, negedge WADDR[8], 1.0);
   $setup(posedge WADDR[9], posedge WCLK, 1.0);
   $setup(negedge WADDR[9], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[9], 1.0);
   $hold(posedge WCLK, negedge WADDR[9], 1.0);
   $setup(posedge WADDR[10], posedge WCLK, 1.0);
   $setup(negedge WADDR[10], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[10], 1.0);
   $hold(posedge WCLK, negedge WADDR[10], 1.0);
   $setup(posedge WDATA[0], posedge WCLK, 1.0);
   $setup(negedge WDATA[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[0], 1.0);
   $hold(posedge WCLK, negedge WDATA[0], 1.0);
   $setup(posedge WDATA[1], posedge WCLK, 1.0);
   $setup(negedge WDATA[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[1], 1.0);
   $hold(posedge WCLK, negedge WDATA[1], 1.0);
   $setup(posedge WDATA[2], posedge WCLK, 1.0);
   $setup(negedge WDATA[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[2], 1.0);
   $hold(posedge WCLK, negedge WDATA[2], 1.0);
   $setup(posedge WDATA[3], posedge WCLK, 1.0);
   $setup(negedge WDATA[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[3], 1.0);
   $hold(posedge WCLK, negedge WDATA[3], 1.0);
   $setup(posedge WDATA[4], posedge WCLK, 1.0);
   $setup(negedge WDATA[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[4], 1.0);
   $hold(posedge WCLK, negedge WDATA[4], 1.0);
   $setup(posedge WDATA[5], posedge WCLK, 1.0);
   $setup(negedge WDATA[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[5], 1.0);
   $hold(posedge WCLK, negedge WDATA[5], 1.0);
   $setup(posedge WDATA[6], posedge WCLK, 1.0);
   $setup(negedge WDATA[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[6], 1.0);
   $hold(posedge WCLK, negedge WDATA[6], 1.0);
   $setup(posedge WDATA[7], posedge WCLK, 1.0);
   $setup(negedge WDATA[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[7], 1.0);
   $hold(posedge WCLK, negedge WDATA[7], 1.0);
   $setup(posedge WCLKE, posedge WCLK, 1.0);
   $setup(negedge WCLKE, posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WCLKE, 1.0);
   $hold(posedge WCLK, negedge WCLKE, 1.0);
   $setup(posedge WE, posedge WCLK, 1.0);
   $setup(negedge WE, posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WE, 1.0);
   $hold(posedge WCLK, negedge WE, 1.0);
   $setup(posedge RADDR[0], posedge RCLKN, 1.0);
   $setup(negedge RADDR[0], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[0], 1.0);
   $hold(posedge RCLKN, negedge RADDR[0], 1.0);
   $setup(posedge RADDR[1], posedge RCLKN, 1.0);
   $setup(negedge RADDR[1], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[1], 1.0);
   $hold(posedge RCLKN, negedge RADDR[1], 1.0);
   $setup(posedge RADDR[2], posedge RCLKN, 1.0);
   $setup(negedge RADDR[2], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[2], 1.0);
   $hold(posedge RCLKN, negedge RADDR[2], 1.0);
   $setup(posedge RADDR[3], posedge RCLKN, 1.0);
   $setup(negedge RADDR[3], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[3], 1.0);
   $hold(posedge RCLKN, negedge RADDR[3], 1.0);
   $setup(posedge RADDR[4], posedge RCLKN, 1.0);
   $setup(negedge RADDR[4], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[4], 1.0);
   $hold(posedge RCLKN, negedge RADDR[4], 1.0);
   $setup(posedge RADDR[5], posedge RCLKN, 1.0);
   $setup(negedge RADDR[5], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[5], 1.0);
   $hold(posedge RCLKN, negedge RADDR[5], 1.0);
   $setup(posedge RADDR[6], posedge RCLKN, 1.0);
   $setup(negedge RADDR[6], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[6], 1.0);
   $hold(posedge RCLKN, negedge RADDR[6], 1.0);
   $setup(posedge RADDR[7], posedge RCLKN, 1.0);
   $setup(negedge RADDR[7], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[7], 1.0);
   $hold(posedge RCLKN, negedge RADDR[7], 1.0);
   $setup(posedge RADDR[8], posedge RCLKN, 1.0);
   $setup(negedge RADDR[8], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[8], 1.0);
   $hold(posedge RCLKN, negedge RADDR[8], 1.0);
   $setup(posedge RADDR[9], posedge RCLKN, 1.0);
   $setup(negedge RADDR[9], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[9], 1.0);
   $hold(posedge RCLKN, negedge RADDR[9], 1.0);
   $setup(posedge RADDR[10], posedge RCLKN, 1.0);
   $setup(negedge RADDR[10], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[10], 1.0);
   $hold(posedge RCLKN, negedge RADDR[10], 1.0);
   $setup(posedge RCLKE, posedge RCLKN, 1.0);
   $setup(negedge RCLKE, posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RCLKE, 1.0);
   $hold(posedge RCLKN, negedge RCLKE, 1.0);
   $setup(posedge RE, posedge RCLKN, 1.0);
   $setup(negedge RE, posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RE, 1.0);
   $hold(posedge RCLKN, negedge RE, 1.0);
endspecify
`endif

endmodule // SB_RAM2048x8NR

//---------------------------------------
//	--- SB_RAM2048x8NW
//---------------------------------------
`timescale 1ps/1ps
module SB_RAM2048x8NW ( RDATA, RCLK, RCLKE, RE, RADDR, WCLKN, WCLKE, WE, WADDR, WDATA ); 

output	[7:0]	RDATA;  
input         	RCLK;   
input           RCLKE; 
input           RE; 
input	[10:0]  RADDR; 
input           WCLKN; 
input           WCLKE; 
input           WE; 
input 	[10:0]  WADDR; 
input 	[7:0]	WDATA; 

parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;


wire WCLK;
assign (weak0, weak1) RCLKE =1'b1 ;
assign (weak0, weak1) RE =1'b0 ;
assign (weak0, weak1) WCLKE =1'b1 ;
assign (weak0, weak1) WE =1'b0 ;
assign WCLK = ~WCLKN;

SB_RAM2048x8  sb_ram2048x8w_inst (
	.RDATA(RDATA),
	.RCLK(RCLK),
	.RCLKE(RCLKE),
	.RE(RE),
	.RADDR(RADDR),
	.WCLK(WCLK),
	.WCLKE(WCLKE),
	.WE(WE),
	.WADDR(WADDR),
	.WDATA(WDATA));

defparam sb_ram2048x8w_inst.INIT_0 = INIT_0;
defparam sb_ram2048x8w_inst.INIT_1 = INIT_1;
defparam sb_ram2048x8w_inst.INIT_2 = INIT_2;
defparam sb_ram2048x8w_inst.INIT_3 = INIT_3;
defparam sb_ram2048x8w_inst.INIT_4 = INIT_4;
defparam sb_ram2048x8w_inst.INIT_5 = INIT_5;
defparam sb_ram2048x8w_inst.INIT_6 = INIT_6;
defparam sb_ram2048x8w_inst.INIT_7 = INIT_7;
defparam sb_ram2048x8w_inst.INIT_8 = INIT_8;
defparam sb_ram2048x8w_inst.INIT_9 = INIT_9;
defparam sb_ram2048x8w_inst.INIT_A = INIT_A;
defparam sb_ram2048x8w_inst.INIT_B = INIT_B;
defparam sb_ram2048x8w_inst.INIT_C = INIT_C;
defparam sb_ram2048x8w_inst.INIT_D = INIT_D;
defparam sb_ram2048x8w_inst.INIT_E = INIT_E;
defparam sb_ram2048x8w_inst.INIT_F = INIT_F;

defparam sb_ram2048x8w_inst.INIT_10 = INIT_10;
defparam sb_ram2048x8w_inst.INIT_11 = INIT_11;
defparam sb_ram2048x8w_inst.INIT_12 = INIT_12;
defparam sb_ram2048x8w_inst.INIT_13 = INIT_13;
defparam sb_ram2048x8w_inst.INIT_14 = INIT_14;
defparam sb_ram2048x8w_inst.INIT_15 = INIT_15;
defparam sb_ram2048x8w_inst.INIT_16 = INIT_16;
defparam sb_ram2048x8w_inst.INIT_17 = INIT_17;
defparam sb_ram2048x8w_inst.INIT_18 = INIT_18;
defparam sb_ram2048x8w_inst.INIT_19 = INIT_19;
defparam sb_ram2048x8w_inst.INIT_1A = INIT_1A;
defparam sb_ram2048x8w_inst.INIT_1B = INIT_1B;
defparam sb_ram2048x8w_inst.INIT_1C = INIT_1C;
defparam sb_ram2048x8w_inst.INIT_1D = INIT_1D;
defparam sb_ram2048x8w_inst.INIT_1E = INIT_1E;
defparam sb_ram2048x8w_inst.INIT_1F = INIT_1F;

defparam sb_ram2048x8w_inst.INIT_20 = INIT_20;
defparam sb_ram2048x8w_inst.INIT_21 = INIT_21;
defparam sb_ram2048x8w_inst.INIT_22 = INIT_22;
defparam sb_ram2048x8w_inst.INIT_23 = INIT_23;
defparam sb_ram2048x8w_inst.INIT_24 = INIT_24;
defparam sb_ram2048x8w_inst.INIT_25 = INIT_25;
defparam sb_ram2048x8w_inst.INIT_26 = INIT_26;
defparam sb_ram2048x8w_inst.INIT_27 = INIT_27;
defparam sb_ram2048x8w_inst.INIT_28 = INIT_28;
defparam sb_ram2048x8w_inst.INIT_29 = INIT_29;
defparam sb_ram2048x8w_inst.INIT_2A = INIT_2A;
defparam sb_ram2048x8w_inst.INIT_2B = INIT_2B;
defparam sb_ram2048x8w_inst.INIT_2C = INIT_2C;
defparam sb_ram2048x8w_inst.INIT_2D = INIT_2D;
defparam sb_ram2048x8w_inst.INIT_2E = INIT_2E;
defparam sb_ram2048x8w_inst.INIT_2F = INIT_2F;

defparam sb_ram2048x8w_inst.INIT_30 = INIT_30;
defparam sb_ram2048x8w_inst.INIT_31 = INIT_31;
defparam sb_ram2048x8w_inst.INIT_32 = INIT_32;
defparam sb_ram2048x8w_inst.INIT_33 = INIT_33;
defparam sb_ram2048x8w_inst.INIT_34 = INIT_34;
defparam sb_ram2048x8w_inst.INIT_35 = INIT_35;
defparam sb_ram2048x8w_inst.INIT_36 = INIT_36;
defparam sb_ram2048x8w_inst.INIT_37 = INIT_37;
defparam sb_ram2048x8w_inst.INIT_38 = INIT_38;
defparam sb_ram2048x8w_inst.INIT_39 = INIT_39;
defparam sb_ram2048x8w_inst.INIT_3A = INIT_3A;
defparam sb_ram2048x8w_inst.INIT_3B = INIT_3B;
defparam sb_ram2048x8w_inst.INIT_3C = INIT_3C;
defparam sb_ram2048x8w_inst.INIT_3D = INIT_3D;
defparam sb_ram2048x8w_inst.INIT_3E = INIT_3E;
defparam sb_ram2048x8w_inst.INIT_3F = INIT_3F;

`ifdef TIMINGCHECK
specify
   (RCLK *> RDATA[0]) = (1.0, 1.0);
   (RCLK *> RDATA[1]) = (1.0, 1.0);
   (RCLK *> RDATA[2]) = (1.0, 1.0);
   (RCLK *> RDATA[3]) = (1.0, 1.0);
   (RCLK *> RDATA[4]) = (1.0, 1.0);
   (RCLK *> RDATA[5]) = (1.0, 1.0);
   (RCLK *> RDATA[6]) = (1.0, 1.0);
   (RCLK *> RDATA[7]) = (1.0, 1.0);
   $setup(posedge WADDR[0], posedge WCLKN, 1.0);
   $setup(negedge WADDR[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[0], 1.0);
   $hold(posedge WCLKN, negedge WADDR[0], 1.0);
   $setup(posedge WADDR[1], posedge WCLKN, 1.0);
   $setup(negedge WADDR[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[1], 1.0);
   $hold(posedge WCLKN, negedge WADDR[1], 1.0);
   $setup(posedge WADDR[2], posedge WCLKN, 1.0);
   $setup(negedge WADDR[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[2], 1.0);
   $hold(posedge WCLKN, negedge WADDR[2], 1.0);
   $setup(posedge WADDR[3], posedge WCLKN, 1.0);
   $setup(negedge WADDR[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[3], 1.0);
   $hold(posedge WCLKN, negedge WADDR[3], 1.0);
   $setup(posedge WADDR[4], posedge WCLKN, 1.0);
   $setup(negedge WADDR[4], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[4], 1.0);
   $hold(posedge WCLKN, negedge WADDR[4], 1.0);
   $setup(posedge WADDR[5], posedge WCLKN, 1.0);
   $setup(negedge WADDR[5], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[5], 1.0);
   $hold(posedge WCLKN, negedge WADDR[5], 1.0);
   $setup(posedge WADDR[6], posedge WCLKN, 1.0);
   $setup(negedge WADDR[6], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[6], 1.0);
   $hold(posedge WCLKN, negedge WADDR[6], 1.0);
   $setup(posedge WADDR[7], posedge WCLKN, 1.0);
   $setup(negedge WADDR[7], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[7], 1.0);
   $hold(posedge WCLKN, negedge WADDR[7], 1.0);
   $setup(posedge WADDR[8], posedge WCLKN, 1.0);
   $setup(negedge WADDR[8], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[8], 1.0);
   $hold(posedge WCLKN, negedge WADDR[8], 1.0);
   $setup(posedge WADDR[9], posedge WCLKN, 1.0);
   $setup(negedge WADDR[9], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[9], 1.0);
   $hold(posedge WCLKN, negedge WADDR[9], 1.0);
   $setup(posedge WADDR[10], posedge WCLKN, 1.0);
   $setup(negedge WADDR[10], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[10], 1.0);
   $hold(posedge WCLKN, negedge WADDR[10], 1.0);
   $setup(posedge WDATA[0], posedge WCLKN, 1.0);
   $setup(negedge WDATA[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[0], 1.0);
   $hold(posedge WCLKN, negedge WDATA[0], 1.0);
   $setup(posedge WDATA[1], posedge WCLKN, 1.0);
   $setup(negedge WDATA[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[1], 1.0);
   $hold(posedge WCLKN, negedge WDATA[1], 1.0);
   $setup(posedge WDATA[2], posedge WCLKN, 1.0);
   $setup(negedge WDATA[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[2], 1.0);
   $hold(posedge WCLKN, negedge WDATA[2], 1.0);
   $setup(posedge WDATA[3], posedge WCLKN, 1.0);
   $setup(negedge WDATA[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[3], 1.0);
   $hold(posedge WCLKN, negedge WDATA[3], 1.0);
   $setup(posedge WDATA[4], posedge WCLKN, 1.0);
   $setup(negedge WDATA[4], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[4], 1.0);
   $hold(posedge WCLKN, negedge WDATA[4], 1.0);
   $setup(posedge WDATA[5], posedge WCLKN, 1.0);
   $setup(negedge WDATA[5], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[5], 1.0);
   $hold(posedge WCLKN, negedge WDATA[5], 1.0);
   $setup(posedge WDATA[6], posedge WCLKN, 1.0);
   $setup(negedge WDATA[6], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[6], 1.0);
   $hold(posedge WCLKN, negedge WDATA[6], 1.0);
   $setup(posedge WDATA[7], posedge WCLKN, 1.0);
   $setup(negedge WDATA[7], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[7], 1.0);
   $hold(posedge WCLKN, negedge WDATA[7], 1.0);
   $setup(posedge WCLKE, posedge WCLKN, 1.0);
   $setup(negedge WCLKE, posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WCLKE, 1.0);
   $hold(posedge WCLKN, negedge WCLKE, 1.0);
   $setup(posedge WE, posedge WCLKN, 1.0);
   $setup(negedge WE, posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WE, 1.0);
   $hold(posedge WCLKN, negedge WE, 1.0);
   $setup(posedge RADDR[0], posedge RCLK, 1.0);
   $setup(negedge RADDR[0], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[0], 1.0);
   $hold(posedge RCLK, negedge RADDR[0], 1.0);
   $setup(posedge RADDR[1], posedge RCLK, 1.0);
   $setup(negedge RADDR[1], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[1], 1.0);
   $hold(posedge RCLK, negedge RADDR[1], 1.0);
   $setup(posedge RADDR[2], posedge RCLK, 1.0);
   $setup(negedge RADDR[2], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[2], 1.0);
   $hold(posedge RCLK, negedge RADDR[2], 1.0);
   $setup(posedge RADDR[3], posedge RCLK, 1.0);
   $setup(negedge RADDR[3], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[3], 1.0);
   $hold(posedge RCLK, negedge RADDR[3], 1.0);
   $setup(posedge RADDR[4], posedge RCLK, 1.0);
   $setup(negedge RADDR[4], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[4], 1.0);
   $hold(posedge RCLK, negedge RADDR[4], 1.0);
   $setup(posedge RADDR[5], posedge RCLK, 1.0);
   $setup(negedge RADDR[5], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[5], 1.0);
   $hold(posedge RCLK, negedge RADDR[5], 1.0);
   $setup(posedge RADDR[6], posedge RCLK, 1.0);
   $setup(negedge RADDR[6], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[6], 1.0);
   $hold(posedge RCLK, negedge RADDR[6], 1.0);
   $setup(posedge RADDR[7], posedge RCLK, 1.0);
   $setup(negedge RADDR[7], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[7], 1.0);
   $hold(posedge RCLK, negedge RADDR[7], 1.0);
   $setup(posedge RADDR[8], posedge RCLK, 1.0);
   $setup(negedge RADDR[8], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[8], 1.0);
   $hold(posedge RCLK, negedge RADDR[8], 1.0);
   $setup(posedge RADDR[9], posedge RCLK, 1.0);
   $setup(negedge RADDR[9], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[9], 1.0);
   $hold(posedge RCLK, negedge RADDR[9], 1.0);
   $setup(posedge RADDR[10], posedge RCLK, 1.0);
   $setup(negedge RADDR[10], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[10], 1.0);
   $hold(posedge RCLK, negedge RADDR[10], 1.0);
   $setup(posedge RCLKE, posedge RCLK, 1.0);
   $setup(negedge RCLKE, posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RCLKE, 1.0);
   $hold(posedge RCLK, negedge RCLKE, 1.0);
   $setup(posedge RE, posedge RCLK, 1.0);
   $setup(negedge RE, posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RE, 1.0);
   $hold(posedge RCLK, negedge RE, 1.0);
endspecify
`endif

endmodule // SB_RAM2048x8NW

//---------------------------------------
//	--- SB_RAM2048x8NRNW
//---------------------------------------
`timescale 1ps/1ps
module SB_RAM2048x8NRNW ( RDATA, RCLKN, RCLKE, RE, RADDR, WCLKN, WCLKE, WE, WADDR, WDATA ); 

output	[7:0]	RDATA;  
input         	RCLKN;   
input           RCLKE; 
input           RE; 
input	[10:0]  RADDR; 
input           WCLKN; 
input           WCLKE; 
input           WE; 
input 	[10:0]  WADDR; 
input 	[7:0]	WDATA;

parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;


wire RCLK, WCLK;
assign (weak0, weak1) RCLKE =1'b1 ;
assign (weak0, weak1) RE =1'b0 ;
assign (weak0, weak1) WCLKE =1'b1 ;
assign (weak0, weak1) WE =1'b0 ;
assign RCLK = ~RCLKN;
assign WCLK = ~WCLKN;

SB_RAM2048x8 sb_ram2048x8rw_inst (
	.RDATA(RDATA),
	.RCLK(RCLK),
	.RCLKE(RCLKE),
	.RE(RE),
	.RADDR(RADDR),
	.WCLK(WCLK),
	.WCLKE(WCLKE),
	.WE(WE),
	.WADDR(WADDR),
	.WDATA(WDATA));

defparam sb_ram2048x8rw_inst.INIT_0 = INIT_0;
defparam sb_ram2048x8rw_inst.INIT_1 = INIT_1;
defparam sb_ram2048x8rw_inst.INIT_2 = INIT_2;
defparam sb_ram2048x8rw_inst.INIT_3 = INIT_3;
defparam sb_ram2048x8rw_inst.INIT_4 = INIT_4;
defparam sb_ram2048x8rw_inst.INIT_5 = INIT_5;
defparam sb_ram2048x8rw_inst.INIT_6 = INIT_6;
defparam sb_ram2048x8rw_inst.INIT_7 = INIT_7;
defparam sb_ram2048x8rw_inst.INIT_8 = INIT_8;
defparam sb_ram2048x8rw_inst.INIT_9 = INIT_9;
defparam sb_ram2048x8rw_inst.INIT_A = INIT_A;
defparam sb_ram2048x8rw_inst.INIT_B = INIT_B;
defparam sb_ram2048x8rw_inst.INIT_C = INIT_C;
defparam sb_ram2048x8rw_inst.INIT_D = INIT_D;
defparam sb_ram2048x8rw_inst.INIT_E = INIT_E;
defparam sb_ram2048x8rw_inst.INIT_F = INIT_F;

defparam sb_ram2048x8rw_inst.INIT_10 = INIT_10;
defparam sb_ram2048x8rw_inst.INIT_11 = INIT_11;
defparam sb_ram2048x8rw_inst.INIT_12 = INIT_12;
defparam sb_ram2048x8rw_inst.INIT_13 = INIT_13;
defparam sb_ram2048x8rw_inst.INIT_14 = INIT_14;
defparam sb_ram2048x8rw_inst.INIT_15 = INIT_15;
defparam sb_ram2048x8rw_inst.INIT_16 = INIT_16;
defparam sb_ram2048x8rw_inst.INIT_17 = INIT_17;
defparam sb_ram2048x8rw_inst.INIT_18 = INIT_18;
defparam sb_ram2048x8rw_inst.INIT_19 = INIT_19;
defparam sb_ram2048x8rw_inst.INIT_1A = INIT_1A;
defparam sb_ram2048x8rw_inst.INIT_1B = INIT_1B;
defparam sb_ram2048x8rw_inst.INIT_1C = INIT_1C;
defparam sb_ram2048x8rw_inst.INIT_1D = INIT_1D;
defparam sb_ram2048x8rw_inst.INIT_1E = INIT_1E;
defparam sb_ram2048x8rw_inst.INIT_1F = INIT_1F;

defparam sb_ram2048x8rw_inst.INIT_20 = INIT_20;
defparam sb_ram2048x8rw_inst.INIT_21 = INIT_21;
defparam sb_ram2048x8rw_inst.INIT_22 = INIT_22;
defparam sb_ram2048x8rw_inst.INIT_23 = INIT_23;
defparam sb_ram2048x8rw_inst.INIT_24 = INIT_24;
defparam sb_ram2048x8rw_inst.INIT_25 = INIT_25;
defparam sb_ram2048x8rw_inst.INIT_26 = INIT_26;
defparam sb_ram2048x8rw_inst.INIT_27 = INIT_27;
defparam sb_ram2048x8rw_inst.INIT_28 = INIT_28;
defparam sb_ram2048x8rw_inst.INIT_29 = INIT_29;
defparam sb_ram2048x8rw_inst.INIT_2A = INIT_2A;
defparam sb_ram2048x8rw_inst.INIT_2B = INIT_2B;
defparam sb_ram2048x8rw_inst.INIT_2C = INIT_2C;
defparam sb_ram2048x8rw_inst.INIT_2D = INIT_2D;
defparam sb_ram2048x8rw_inst.INIT_2E = INIT_2E;
defparam sb_ram2048x8rw_inst.INIT_2F = INIT_2F;

defparam sb_ram2048x8rw_inst.INIT_30 = INIT_30;
defparam sb_ram2048x8rw_inst.INIT_31 = INIT_31;
defparam sb_ram2048x8rw_inst.INIT_32 = INIT_32;
defparam sb_ram2048x8rw_inst.INIT_33 = INIT_33;
defparam sb_ram2048x8rw_inst.INIT_34 = INIT_34;
defparam sb_ram2048x8rw_inst.INIT_35 = INIT_35;
defparam sb_ram2048x8rw_inst.INIT_36 = INIT_36;
defparam sb_ram2048x8rw_inst.INIT_37 = INIT_37;
defparam sb_ram2048x8rw_inst.INIT_38 = INIT_38;
defparam sb_ram2048x8rw_inst.INIT_39 = INIT_39;
defparam sb_ram2048x8rw_inst.INIT_3A = INIT_3A;
defparam sb_ram2048x8rw_inst.INIT_3B = INIT_3B;
defparam sb_ram2048x8rw_inst.INIT_3C = INIT_3C;
defparam sb_ram2048x8rw_inst.INIT_3D = INIT_3D;
defparam sb_ram2048x8rw_inst.INIT_3E = INIT_3E;
defparam sb_ram2048x8rw_inst.INIT_3F = INIT_3F;

`ifdef TIMINGCHECK
specify
   (RCLKN *> RDATA[0]) = (1.0, 1.0);
   (RCLKN *> RDATA[1]) = (1.0, 1.0);
   (RCLKN *> RDATA[2]) = (1.0, 1.0);
   (RCLKN *> RDATA[3]) = (1.0, 1.0);
   (RCLKN *> RDATA[4]) = (1.0, 1.0);
   (RCLKN *> RDATA[5]) = (1.0, 1.0);
   (RCLKN *> RDATA[6]) = (1.0, 1.0);
   (RCLKN *> RDATA[7]) = (1.0, 1.0);
   $setup(posedge WADDR[0], posedge WCLKN, 1.0);
   $setup(negedge WADDR[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[0], 1.0);
   $hold(posedge WCLKN, negedge WADDR[0], 1.0);
   $setup(posedge WADDR[1], posedge WCLKN, 1.0);
   $setup(negedge WADDR[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[1], 1.0);
   $hold(posedge WCLKN, negedge WADDR[1], 1.0);
   $setup(posedge WADDR[2], posedge WCLKN, 1.0);
   $setup(negedge WADDR[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[2], 1.0);
   $hold(posedge WCLKN, negedge WADDR[2], 1.0);
   $setup(posedge WADDR[3], posedge WCLKN, 1.0);
   $setup(negedge WADDR[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[3], 1.0);
   $hold(posedge WCLKN, negedge WADDR[3], 1.0);
   $setup(posedge WADDR[4], posedge WCLKN, 1.0);
   $setup(negedge WADDR[4], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[4], 1.0);
   $hold(posedge WCLKN, negedge WADDR[4], 1.0);
   $setup(posedge WADDR[5], posedge WCLKN, 1.0);
   $setup(negedge WADDR[5], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[5], 1.0);
   $hold(posedge WCLKN, negedge WADDR[5], 1.0);
   $setup(posedge WADDR[6], posedge WCLKN, 1.0);
   $setup(negedge WADDR[6], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[6], 1.0);
   $hold(posedge WCLKN, negedge WADDR[6], 1.0);
   $setup(posedge WADDR[7], posedge WCLKN, 1.0);
   $setup(negedge WADDR[7], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[7], 1.0);
   $hold(posedge WCLKN, negedge WADDR[7], 1.0);
   $setup(posedge WADDR[8], posedge WCLKN, 1.0);
   $setup(negedge WADDR[8], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[8], 1.0);
   $hold(posedge WCLKN, negedge WADDR[8], 1.0);
   $setup(posedge WADDR[9], posedge WCLKN, 1.0);
   $setup(negedge WADDR[9], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[9], 1.0);
   $hold(posedge WCLKN, negedge WADDR[9], 1.0);
   $setup(posedge WADDR[10], posedge WCLKN, 1.0);
   $setup(negedge WADDR[10], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[10], 1.0);
   $hold(posedge WCLKN, negedge WADDR[10], 1.0);
   $setup(posedge WDATA[0], posedge WCLKN, 1.0);
   $setup(negedge WDATA[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[0], 1.0);
   $hold(posedge WCLKN, negedge WDATA[0], 1.0);
   $setup(posedge WDATA[1], posedge WCLKN, 1.0);
   $setup(negedge WDATA[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[1], 1.0);
   $hold(posedge WCLKN, negedge WDATA[1], 1.0);
   $setup(posedge WDATA[2], posedge WCLKN, 1.0);
   $setup(negedge WDATA[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[2], 1.0);
   $hold(posedge WCLKN, negedge WDATA[2], 1.0);
   $setup(posedge WDATA[3], posedge WCLKN, 1.0);
   $setup(negedge WDATA[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[3], 1.0);
   $hold(posedge WCLKN, negedge WDATA[3], 1.0);
   $setup(posedge WDATA[4], posedge WCLKN, 1.0);
   $setup(negedge WDATA[4], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[4], 1.0);
   $hold(posedge WCLKN, negedge WDATA[4], 1.0);
   $setup(posedge WDATA[5], posedge WCLKN, 1.0);
   $setup(negedge WDATA[5], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[5], 1.0);
   $hold(posedge WCLKN, negedge WDATA[5], 1.0);
   $setup(posedge WDATA[6], posedge WCLKN, 1.0);
   $setup(negedge WDATA[6], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[6], 1.0);
   $hold(posedge WCLKN, negedge WDATA[6], 1.0);
   $setup(posedge WDATA[7], posedge WCLKN, 1.0);
   $setup(negedge WDATA[7], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[7], 1.0);
   $hold(posedge WCLKN, negedge WDATA[7], 1.0);
   $setup(posedge WCLKE, posedge WCLKN, 1.0);
   $setup(negedge WCLKE, posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WCLKE, 1.0);
   $hold(posedge WCLKN, negedge WCLKE, 1.0);
   $setup(posedge WE, posedge WCLKN, 1.0);
   $setup(negedge WE, posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WE, 1.0);
   $hold(posedge WCLKN, negedge WE, 1.0);
   $setup(posedge RADDR[0], posedge RCLKN, 1.0);
   $setup(negedge RADDR[0], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[0], 1.0);
   $hold(posedge RCLKN, negedge RADDR[0], 1.0);
   $setup(posedge RADDR[1], posedge RCLKN, 1.0);
   $setup(negedge RADDR[1], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[1], 1.0);
   $hold(posedge RCLKN, negedge RADDR[1], 1.0);
   $setup(posedge RADDR[2], posedge RCLKN, 1.0);
   $setup(negedge RADDR[2], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[2], 1.0);
   $hold(posedge RCLKN, negedge RADDR[2], 1.0);
   $setup(posedge RADDR[3], posedge RCLKN, 1.0);
   $setup(negedge RADDR[3], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[3], 1.0);
   $hold(posedge RCLKN, negedge RADDR[3], 1.0);
   $setup(posedge RADDR[4], posedge RCLKN, 1.0);
   $setup(negedge RADDR[4], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[4], 1.0);
   $hold(posedge RCLKN, negedge RADDR[4], 1.0);
   $setup(posedge RADDR[5], posedge RCLKN, 1.0);
   $setup(negedge RADDR[5], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[5], 1.0);
   $hold(posedge RCLKN, negedge RADDR[5], 1.0);
   $setup(posedge RADDR[6], posedge RCLKN, 1.0);
   $setup(negedge RADDR[6], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[6], 1.0);
   $hold(posedge RCLKN, negedge RADDR[6], 1.0);
   $setup(posedge RADDR[7], posedge RCLKN, 1.0);
   $setup(negedge RADDR[7], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[7], 1.0);
   $hold(posedge RCLKN, negedge RADDR[7], 1.0);
   $setup(posedge RADDR[8], posedge RCLKN, 1.0);
   $setup(negedge RADDR[8], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[8], 1.0);
   $hold(posedge RCLKN, negedge RADDR[8], 1.0);
   $setup(posedge RADDR[9], posedge RCLKN, 1.0);
   $setup(negedge RADDR[9], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[9], 1.0);
   $hold(posedge RCLKN, negedge RADDR[9], 1.0);
   $setup(posedge RADDR[10], posedge RCLKN, 1.0);
   $setup(negedge RADDR[10], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[10], 1.0);
   $hold(posedge RCLKN, negedge RADDR[10], 1.0);
   $setup(posedge RCLKE, posedge RCLKN, 1.0);
   $setup(negedge RCLKE, posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RCLKE, 1.0);
   $hold(posedge RCLKN, negedge RCLKE, 1.0);
   $setup(posedge RE, posedge RCLKN, 1.0);
   $setup(negedge RE, posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RE, 1.0);
   $hold(posedge RCLKN, negedge RE, 1.0);
endspecify
`endif

endmodule // SB_RAM2048x8NRNW 

//---------------------------------------
//	--- SB_RAM4096x4
//---------------------------------------
`timescale 1ps/1ps
module SB_RAM4096x4 ( RDATA, RCLK, RCLKE, RE, RADDR, WCLK, WCLKE, WE, WADDR, WDATA ); 

output	[3:0]	RDATA;  
input         	RCLK;   
input           RCLKE; 
input           RE; 
input	[11:0]  RADDR; 
input           WCLK; 
input           WCLKE; 
input           WE; 
input 	[11:0]  WADDR; 
input 	[3:0]	WDATA;

parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

// local Parameters
localparam			CLOCK_PERIOD = 200;	//
localparam 			DELAY	= (CLOCK_PERIOD/10);		// Clock-to-output delay. Zero
							// time delays can be confusing
							// and sometimes cause problems.
localparam 			BUS_WIDTH = 4;		// Width of RAM (number of bits)

localparam 			ADDRESS_BUS_SIZE = 12;	// Number of bits required to
							// represent the RAM address

localparam   ADDRESSABLE_SPACE  = 2**ADDRESS_BUS_SIZE;	// Decimal address range [2^Size:0]


// SIGNAL DECLARATIONS
wire			   	WCLK_g, RCLK_g;
reg 				WCLKE_sync, RCLKE_sync; 
assign (weak0, weak1) RCLKE =1'b1 ;
assign (weak0, weak1) RE =1'b0 ;
assign (weak0, weak1) WCLKE =1'b1 ;
assign (weak0, weak1) WE =1'b0 ;
reg	Memory	[BUS_WIDTH*ADDRESSABLE_SPACE-1:0];
// 
event Read_e, Write_e;

//////////////////// Collision detect begins here ///////////////////////////////
localparam 	TRUE = 1'b1;
localparam	FALSE = 1'b0;
reg 		Time_Collision_Detected = 1'b0;
wire		Address_Collision_Detected;

event Collision_e;

time COLLISION_TIME_WINDOW = (CLOCK_PERIOD/8); // This is an arbitray value, but is better than using an absolute 
						    // value, because the actual time window depends on the actual silicon 
						    // implementation. Thus the test is indicative of an Error and not
						    // guaranteed to be an error. Even so this is usefull.
time time_WCLK_RCLK, time_WCLK, time_RCLK;


//function reg Check_Timed_Window_Violation;
function	Check_Timed_Window_Violation;	
input T1, T2, Minimum_Time_Window;
time T1, T2;
time Minimum_Time_Window;
time Difference;	
	begin
		Difference = (T1 - T2);
		if (Difference < 0) Difference = -Difference;
		Check_Timed_Window_Violation = (Difference < Minimum_Time_Window);
	end
endfunction


initial begin
       time_WCLK = CLOCK_PERIOD;	// Arbitrary initialisation value, ensure no window collison error on first clock edge.
       time_RCLK = (CLOCK_PERIOD*8);	// Arbitrary initialisation difference value, ensure no collision error on first clock edge.					
end

integer	i,j;


initial	//	initialize ram_16k (4096x4) by init parameters, section by section
begin
	for	(i=0; i<=(256/BUS_WIDTH)-1; i=i+1)       
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)    
		begin 

			Memory[BUS_WIDTH*i+j]		=	INIT_0[BUS_WIDTH*i+j];
			Memory[256*1+BUS_WIDTH*i+j]	=	INIT_1[BUS_WIDTH*i+j];
			Memory[256*2+BUS_WIDTH*i+j]	=	INIT_2[BUS_WIDTH*i+j];
			Memory[256*3+BUS_WIDTH*i+j]	=	INIT_3[BUS_WIDTH*i+j];
			Memory[256*4+BUS_WIDTH*i+j]	=	INIT_4[BUS_WIDTH*i+j];
			Memory[256*5+BUS_WIDTH*i+j]	=	INIT_5[BUS_WIDTH*i+j];
			Memory[256*6+BUS_WIDTH*i+j]	=	INIT_6[BUS_WIDTH*i+j];
			Memory[256*7+BUS_WIDTH*i+j]	=	INIT_7[BUS_WIDTH*i+j];
			Memory[256*8+BUS_WIDTH*i+j]	=	INIT_8[BUS_WIDTH*i+j];
			Memory[256*9+BUS_WIDTH*i+j]	=	INIT_9[BUS_WIDTH*i+j];
			Memory[256*10+BUS_WIDTH*i+j]	=	INIT_A[BUS_WIDTH*i+j];
			Memory[256*11+BUS_WIDTH*i+j]	=	INIT_B[BUS_WIDTH*i+j];
			Memory[256*12+BUS_WIDTH*i+j]	=	INIT_C[BUS_WIDTH*i+j];
			Memory[256*13+BUS_WIDTH*i+j]	=	INIT_D[BUS_WIDTH*i+j];
			Memory[256*14+BUS_WIDTH*i+j]	=	INIT_E[BUS_WIDTH*i+j];
			Memory[256*15+BUS_WIDTH*i+j]	=	INIT_F[BUS_WIDTH*i+j];

			Memory[256*16+BUS_WIDTH*i+j]	=	INIT_10[BUS_WIDTH*i+j];
			Memory[256*17+BUS_WIDTH*i+j]	=	INIT_11[BUS_WIDTH*i+j];
			Memory[256*18+BUS_WIDTH*i+j]	=	INIT_12[BUS_WIDTH*i+j];
			Memory[256*19+BUS_WIDTH*i+j]	=	INIT_13[BUS_WIDTH*i+j];
			Memory[256*20+BUS_WIDTH*i+j]	=	INIT_14[BUS_WIDTH*i+j];
			Memory[256*21+BUS_WIDTH*i+j]	=	INIT_15[BUS_WIDTH*i+j];
			Memory[256*22+BUS_WIDTH*i+j]	=	INIT_16[BUS_WIDTH*i+j];
			Memory[256*23+BUS_WIDTH*i+j]	=	INIT_17[BUS_WIDTH*i+j];
			Memory[256*24+BUS_WIDTH*i+j]	=	INIT_18[BUS_WIDTH*i+j];
			Memory[256*25+BUS_WIDTH*i+j]	=	INIT_19[BUS_WIDTH*i+j];
			Memory[256*26+BUS_WIDTH*i+j]	=	INIT_1A[BUS_WIDTH*i+j];
			Memory[256*27+BUS_WIDTH*i+j]	=	INIT_1B[BUS_WIDTH*i+j];
			Memory[256*28+BUS_WIDTH*i+j]	=	INIT_1C[BUS_WIDTH*i+j];
			Memory[256*29+BUS_WIDTH*i+j]	=	INIT_1D[BUS_WIDTH*i+j];
			Memory[256*30+BUS_WIDTH*i+j]	=	INIT_1E[BUS_WIDTH*i+j];
			Memory[256*31+BUS_WIDTH*i+j]	=	INIT_1F[BUS_WIDTH*i+j];

			Memory[256*32+BUS_WIDTH*i+j]	=	INIT_20[BUS_WIDTH*i+j];
			Memory[256*33+BUS_WIDTH*i+j]	=	INIT_21[BUS_WIDTH*i+j];
			Memory[256*34+BUS_WIDTH*i+j]	=	INIT_22[BUS_WIDTH*i+j];
			Memory[256*35+BUS_WIDTH*i+j]	=	INIT_23[BUS_WIDTH*i+j];
			Memory[256*36+BUS_WIDTH*i+j]	=	INIT_24[BUS_WIDTH*i+j];
			Memory[256*37+BUS_WIDTH*i+j]	=	INIT_25[BUS_WIDTH*i+j];
			Memory[256*38+BUS_WIDTH*i+j]	=	INIT_26[BUS_WIDTH*i+j];
			Memory[256*39+BUS_WIDTH*i+j]	=	INIT_27[BUS_WIDTH*i+j];
			Memory[256*40+BUS_WIDTH*i+j]	=	INIT_28[BUS_WIDTH*i+j];
			Memory[256*41+BUS_WIDTH*i+j]	=	INIT_29[BUS_WIDTH*i+j];
			Memory[256*42+BUS_WIDTH*i+j]	=	INIT_2A[BUS_WIDTH*i+j];
			Memory[256*43+BUS_WIDTH*i+j]	=	INIT_2B[BUS_WIDTH*i+j];
			Memory[256*44+BUS_WIDTH*i+j]	=	INIT_2C[BUS_WIDTH*i+j];
			Memory[256*45+BUS_WIDTH*i+j]	=	INIT_2D[BUS_WIDTH*i+j];
			Memory[256*46+BUS_WIDTH*i+j]	=	INIT_2E[BUS_WIDTH*i+j];
			Memory[256*47+BUS_WIDTH*i+j]	=	INIT_2F[BUS_WIDTH*i+j];

			Memory[256*48+BUS_WIDTH*i+j]	=	INIT_30[BUS_WIDTH*i+j];
			Memory[256*49+BUS_WIDTH*i+j]	=	INIT_31[BUS_WIDTH*i+j];
			Memory[256*50+BUS_WIDTH*i+j]	=	INIT_32[BUS_WIDTH*i+j];
			Memory[256*51+BUS_WIDTH*i+j]	=	INIT_33[BUS_WIDTH*i+j];
			Memory[256*52+BUS_WIDTH*i+j]	=	INIT_34[BUS_WIDTH*i+j];
			Memory[256*53+BUS_WIDTH*i+j]	=	INIT_35[BUS_WIDTH*i+j];
			Memory[256*54+BUS_WIDTH*i+j]	=	INIT_36[BUS_WIDTH*i+j];
			Memory[256*55+BUS_WIDTH*i+j]	=	INIT_37[BUS_WIDTH*i+j];
			Memory[256*56+BUS_WIDTH*i+j]	=	INIT_38[BUS_WIDTH*i+j];
			Memory[256*57+BUS_WIDTH*i+j]	=	INIT_39[BUS_WIDTH*i+j];
			Memory[256*58+BUS_WIDTH*i+j]	=	INIT_3A[BUS_WIDTH*i+j];
			Memory[256*59+BUS_WIDTH*i+j]	=	INIT_3B[BUS_WIDTH*i+j];
			Memory[256*60+BUS_WIDTH*i+j]	=	INIT_3C[BUS_WIDTH*i+j];
			Memory[256*61+BUS_WIDTH*i+j]	=	INIT_3D[BUS_WIDTH*i+j];
			Memory[256*62+BUS_WIDTH*i+j]	=	INIT_3E[BUS_WIDTH*i+j];
			Memory[256*63+BUS_WIDTH*i+j]	=	INIT_3F[BUS_WIDTH*i+j];

		end 
	end

end

assign Address_Collision_Detected = ((RE & WE & WCLKE & RCLKE)&(WADDR == RADDR)); 

always @(WCLK or WCLKE) 
begin 
	if(~WCLK)
	WCLKE_sync = WCLKE;   	
end 

always @(RCLK or RCLKE) 
begin 
	if (~RCLK)
	RCLKE_sync = RCLKE; 	
end 

assign WCLK_g = WCLK & WCLKE_sync;
assign RCLK_g = RCLK & RCLKE_sync;


always @(posedge WCLK_g) begin
	time_WCLK = $time;
end

always @(posedge RCLK_g) begin
    	time_RCLK = $time;
end
integer	SB_RAM4096x4_RDATA_log_file;					//.....................
initial	SB_RAM4096x4_RDATA_log_file=("SB_RAM4096x4_RDATA_log_file.txt");	//.....................
always @(posedge WCLK_g) begin

	Time_Collision_Detected = Check_Timed_Window_Violation(time_WCLK,time_RCLK,COLLISION_TIME_WINDOW);
        if (Time_Collision_Detected & Address_Collision_Detected)begin
        	$display("Warning: Write-Read collision detected, Data read value is XXXX\n");
 		$display("WCLK Time: %.3f   RCLK Time:%.3f  ",time_WCLK, time_RCLK,"WADDR: %d   RADDR:%d\n",WADDR, RADDR); 
 		$fdisplay(SB_RAM4096x4_RDATA_log_file,"Warning: Write-Read collision detected, Data read value is XXXX\n");
		$fdisplay(SB_RAM4096x4_RDATA_log_file,"WCLK Time: %.3f   RCLK Time:%.3f  ",time_WCLK, time_RCLK, "WADDR: %d   RADDR:%d\n",WADDR, RADDR); 	
 		-> Collision_e;
	end
end

//	code modify for universal verilog compiler

always @ (posedge WCLK_g)
begin
	if	(WE)
	begin
		-> Write_e;
		for	(i=0;i<=BUS_WIDTH-1; i=i+1)
		begin
				Memory[WADDR*BUS_WIDTH+i]	<=	WDATA[i];
		end
	end
end

reg	[BUS_WIDTH-1:0]	RDATA = 0;

// Look at the rising edge of the clock

always @ (posedge RCLK_g)
begin
	if	(RE)
	begin
		-> Read_e;
		if	(Time_Collision_Detected & Address_Collision_Detected) 
			RDATA <= 16'hXXXX;
		else
			for	(i=0;i<=BUS_WIDTH-1;i=i+1)
				RDATA[i]	<= Memory[RADDR*BUS_WIDTH+i];
	end
end

`ifdef TIMINGCHECK
specify
   (RCLK *> RDATA[0]) = (1.0, 1.0);
   (RCLK *> RDATA[1]) = (1.0, 1.0);
   (RCLK *> RDATA[2]) = (1.0, 1.0);
   (RCLK *> RDATA[3]) = (1.0, 1.0);
   $setup(posedge WADDR[0], posedge WCLK, 1.0);
   $setup(negedge WADDR[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[0], 1.0);
   $hold(posedge WCLK, negedge WADDR[0], 1.0);
   $setup(posedge WADDR[1], posedge WCLK, 1.0);
   $setup(negedge WADDR[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[1], 1.0);
   $hold(posedge WCLK, negedge WADDR[1], 1.0);
   $setup(posedge WADDR[2], posedge WCLK, 1.0);
   $setup(negedge WADDR[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[2], 1.0);
   $hold(posedge WCLK, negedge WADDR[2], 1.0);
   $setup(posedge WADDR[3], posedge WCLK, 1.0);
   $setup(negedge WADDR[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[3], 1.0);
   $hold(posedge WCLK, negedge WADDR[3], 1.0);
   $setup(posedge WADDR[4], posedge WCLK, 1.0);
   $setup(negedge WADDR[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[4], 1.0);
   $hold(posedge WCLK, negedge WADDR[4], 1.0);
   $setup(posedge WADDR[5], posedge WCLK, 1.0);
   $setup(negedge WADDR[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[5], 1.0);
   $hold(posedge WCLK, negedge WADDR[5], 1.0);
   $setup(posedge WADDR[6], posedge WCLK, 1.0);
   $setup(negedge WADDR[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[6], 1.0);
   $hold(posedge WCLK, negedge WADDR[6], 1.0);
   $setup(posedge WADDR[7], posedge WCLK, 1.0);
   $setup(negedge WADDR[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[7], 1.0);
   $hold(posedge WCLK, negedge WADDR[7], 1.0);
   $setup(posedge WADDR[8], posedge WCLK, 1.0);
   $setup(negedge WADDR[8], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[8], 1.0);
   $hold(posedge WCLK, negedge WADDR[8], 1.0);
   $setup(posedge WADDR[9], posedge WCLK, 1.0);
   $setup(negedge WADDR[9], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[9], 1.0);
   $hold(posedge WCLK, negedge WADDR[9], 1.0);
   $setup(posedge WADDR[10], posedge WCLK, 1.0);
   $setup(negedge WADDR[10], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[10], 1.0);
   $hold(posedge WCLK, negedge WADDR[10], 1.0);
   $setup(posedge WADDR[11], posedge WCLK, 1.0);
   $setup(negedge WADDR[11], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[11], 1.0);
   $hold(posedge WCLK, negedge WADDR[11], 1.0);
   $setup(posedge WDATA[0], posedge WCLK, 1.0);
   $setup(negedge WDATA[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[0], 1.0);
   $hold(posedge WCLK, negedge WDATA[0], 1.0);
   $setup(posedge WDATA[1], posedge WCLK, 1.0);
   $setup(negedge WDATA[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[1], 1.0);
   $hold(posedge WCLK, negedge WDATA[1], 1.0);
   $setup(posedge WDATA[2], posedge WCLK, 1.0);
   $setup(negedge WDATA[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[2], 1.0);
   $hold(posedge WCLK, negedge WDATA[2], 1.0);
   $setup(posedge WDATA[3], posedge WCLK, 1.0);
   $setup(negedge WDATA[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[3], 1.0);
   $hold(posedge WCLK, negedge WDATA[3], 1.0);
   $setup(posedge WCLKE, posedge WCLK, 1.0);
   $setup(negedge WCLKE, posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WCLKE, 1.0);
   $hold(posedge WCLK, negedge WCLKE, 1.0);
   $setup(posedge WE, posedge WCLK, 1.0);
   $setup(negedge WE, posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WE, 1.0);
   $hold(posedge WCLK, negedge WE, 1.0);
   $setup(posedge RADDR[0], posedge RCLK, 1.0);
   $setup(negedge RADDR[0], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[0], 1.0);
   $hold(posedge RCLK, negedge RADDR[0], 1.0);
   $setup(posedge RADDR[1], posedge RCLK, 1.0);
   $setup(negedge RADDR[1], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[1], 1.0);
   $hold(posedge RCLK, negedge RADDR[1], 1.0);
   $setup(posedge RADDR[2], posedge RCLK, 1.0);
   $setup(negedge RADDR[2], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[2], 1.0);
   $hold(posedge RCLK, negedge RADDR[2], 1.0);
   $setup(posedge RADDR[3], posedge RCLK, 1.0);
   $setup(negedge RADDR[3], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[3], 1.0);
   $hold(posedge RCLK, negedge RADDR[3], 1.0);
   $setup(posedge RADDR[4], posedge RCLK, 1.0);
   $setup(negedge RADDR[4], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[4], 1.0);
   $hold(posedge RCLK, negedge RADDR[4], 1.0);
   $setup(posedge RADDR[5], posedge RCLK, 1.0);
   $setup(negedge RADDR[5], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[5], 1.0);
   $hold(posedge RCLK, negedge RADDR[5], 1.0);
   $setup(posedge RADDR[6], posedge RCLK, 1.0);
   $setup(negedge RADDR[6], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[6], 1.0);
   $hold(posedge RCLK, negedge RADDR[6], 1.0);
   $setup(posedge RADDR[7], posedge RCLK, 1.0);
   $setup(negedge RADDR[7], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[7], 1.0);
   $hold(posedge RCLK, negedge RADDR[7], 1.0);
   $setup(posedge RADDR[8], posedge RCLK, 1.0);
   $setup(negedge RADDR[8], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[8], 1.0);
   $hold(posedge RCLK, negedge RADDR[8], 1.0);
   $setup(posedge RADDR[9], posedge RCLK, 1.0);
   $setup(negedge RADDR[9], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[9], 1.0);
   $hold(posedge RCLK, negedge RADDR[9], 1.0);
   $setup(posedge RADDR[10], posedge RCLK, 1.0);
   $setup(negedge RADDR[10], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[10], 1.0);
   $hold(posedge RCLK, negedge RADDR[10], 1.0);
   $setup(posedge RADDR[11], posedge RCLK, 1.0);
   $setup(negedge RADDR[11], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[11], 1.0);
   $hold(posedge RCLK, negedge RADDR[11], 1.0);
   $setup(posedge RCLKE, posedge RCLK, 1.0);
   $setup(negedge RCLKE, posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RCLKE, 1.0);
   $hold(posedge RCLK, negedge RCLKE, 1.0);
   $setup(posedge RE, posedge RCLK, 1.0);
   $setup(negedge RE, posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RE, 1.0);
   $hold(posedge RCLK, negedge RE, 1.0);
endspecify
`endif

endmodule // SB_RAM4096x4

//---------------------------------------
//	--- SB_RAM4096x4NR
//---------------------------------------
`timescale 1ps/1ps
module SB_RAM4096x4NR ( RDATA, RCLKN, RCLKE, RE, RADDR, WCLK, WCLKE, WE, WADDR, WDATA ); 

output	[3:0]	RDATA;  
input         	RCLKN;   
input           RCLKE; 
input           RE; 
input	[11:0]  RADDR; 
input           WCLK; 
input           WCLKE; 
input           WE; 
input 	[11:0]  WADDR; 
input 	[3:0]	WDATA; 
 
parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;


wire RCLK;
assign (weak0, weak1) RCLKE =1'b1 ;
assign (weak0, weak1) RE =1'b0 ;
assign (weak0, weak1) WCLKE =1'b1 ;
assign (weak0, weak1) WE =1'b0 ;
assign RCLK = ~RCLKN;

SB_RAM4096x4 sb_ram4096x4r_inst (
	.RDATA(RDATA),
	.RCLK(RCLK),
	.RCLKE(RCLKE),
	.RE(RE),
	.RADDR(RADDR),
	.WCLK(WCLK),
	.WCLKE(WCLKE),
	.WE(WE),
	.WADDR(WADDR),
	.WDATA(WDATA));

defparam sb_ram4096x4r_inst.INIT_0 = INIT_0;
defparam sb_ram4096x4r_inst.INIT_1 = INIT_1;
defparam sb_ram4096x4r_inst.INIT_2 = INIT_2;
defparam sb_ram4096x4r_inst.INIT_3 = INIT_3;
defparam sb_ram4096x4r_inst.INIT_4 = INIT_4;
defparam sb_ram4096x4r_inst.INIT_5 = INIT_5;
defparam sb_ram4096x4r_inst.INIT_6 = INIT_6;
defparam sb_ram4096x4r_inst.INIT_7 = INIT_7;
defparam sb_ram4096x4r_inst.INIT_8 = INIT_8;
defparam sb_ram4096x4r_inst.INIT_9 = INIT_9;
defparam sb_ram4096x4r_inst.INIT_A = INIT_A;
defparam sb_ram4096x4r_inst.INIT_B = INIT_B;
defparam sb_ram4096x4r_inst.INIT_C = INIT_C;
defparam sb_ram4096x4r_inst.INIT_D = INIT_D;
defparam sb_ram4096x4r_inst.INIT_E = INIT_E;
defparam sb_ram4096x4r_inst.INIT_F = INIT_F;

defparam sb_ram4096x4r_inst.INIT_10 = INIT_10;
defparam sb_ram4096x4r_inst.INIT_11 = INIT_11;
defparam sb_ram4096x4r_inst.INIT_12 = INIT_12;
defparam sb_ram4096x4r_inst.INIT_13 = INIT_13;
defparam sb_ram4096x4r_inst.INIT_14 = INIT_14;
defparam sb_ram4096x4r_inst.INIT_15 = INIT_15;
defparam sb_ram4096x4r_inst.INIT_16 = INIT_16;
defparam sb_ram4096x4r_inst.INIT_17 = INIT_17;
defparam sb_ram4096x4r_inst.INIT_18 = INIT_18;
defparam sb_ram4096x4r_inst.INIT_19 = INIT_19;
defparam sb_ram4096x4r_inst.INIT_1A = INIT_1A;
defparam sb_ram4096x4r_inst.INIT_1B = INIT_1B;
defparam sb_ram4096x4r_inst.INIT_1C = INIT_1C;
defparam sb_ram4096x4r_inst.INIT_1D = INIT_1D;
defparam sb_ram4096x4r_inst.INIT_1E = INIT_1E;
defparam sb_ram4096x4r_inst.INIT_1F = INIT_1F;

defparam sb_ram4096x4r_inst.INIT_20 = INIT_20;
defparam sb_ram4096x4r_inst.INIT_21 = INIT_21;
defparam sb_ram4096x4r_inst.INIT_22 = INIT_22;
defparam sb_ram4096x4r_inst.INIT_23 = INIT_23;
defparam sb_ram4096x4r_inst.INIT_24 = INIT_24;
defparam sb_ram4096x4r_inst.INIT_25 = INIT_25;
defparam sb_ram4096x4r_inst.INIT_26 = INIT_26;
defparam sb_ram4096x4r_inst.INIT_27 = INIT_27;
defparam sb_ram4096x4r_inst.INIT_28 = INIT_28;
defparam sb_ram4096x4r_inst.INIT_29 = INIT_29;
defparam sb_ram4096x4r_inst.INIT_2A = INIT_2A;
defparam sb_ram4096x4r_inst.INIT_2B = INIT_2B;
defparam sb_ram4096x4r_inst.INIT_2C = INIT_2C;
defparam sb_ram4096x4r_inst.INIT_2D = INIT_2D;
defparam sb_ram4096x4r_inst.INIT_2E = INIT_2E;
defparam sb_ram4096x4r_inst.INIT_2F = INIT_2F;

defparam sb_ram4096x4r_inst.INIT_30 = INIT_30;
defparam sb_ram4096x4r_inst.INIT_31 = INIT_31;
defparam sb_ram4096x4r_inst.INIT_32 = INIT_32;
defparam sb_ram4096x4r_inst.INIT_33 = INIT_33;
defparam sb_ram4096x4r_inst.INIT_34 = INIT_34;
defparam sb_ram4096x4r_inst.INIT_35 = INIT_35;
defparam sb_ram4096x4r_inst.INIT_36 = INIT_36;
defparam sb_ram4096x4r_inst.INIT_37 = INIT_37;
defparam sb_ram4096x4r_inst.INIT_38 = INIT_38;
defparam sb_ram4096x4r_inst.INIT_39 = INIT_39;
defparam sb_ram4096x4r_inst.INIT_3A = INIT_3A;
defparam sb_ram4096x4r_inst.INIT_3B = INIT_3B;
defparam sb_ram4096x4r_inst.INIT_3C = INIT_3C;
defparam sb_ram4096x4r_inst.INIT_3D = INIT_3D;
defparam sb_ram4096x4r_inst.INIT_3E = INIT_3E;
defparam sb_ram4096x4r_inst.INIT_3F = INIT_3F;


`ifdef TIMINGCHECK
specify
   (RCLKN *> RDATA[0]) = (1.0, 1.0);
   (RCLKN *> RDATA[1]) = (1.0, 1.0);
   (RCLKN *> RDATA[2]) = (1.0, 1.0);
   (RCLKN *> RDATA[3]) = (1.0, 1.0);
   $setup(posedge WADDR[0], posedge WCLK, 1.0);
   $setup(negedge WADDR[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[0], 1.0);
   $hold(posedge WCLK, negedge WADDR[0], 1.0);
   $setup(posedge WADDR[1], posedge WCLK, 1.0);
   $setup(negedge WADDR[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[1], 1.0);
   $hold(posedge WCLK, negedge WADDR[1], 1.0);
   $setup(posedge WADDR[2], posedge WCLK, 1.0);
   $setup(negedge WADDR[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[2], 1.0);
   $hold(posedge WCLK, negedge WADDR[2], 1.0);
   $setup(posedge WADDR[3], posedge WCLK, 1.0);
   $setup(negedge WADDR[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[3], 1.0);
   $hold(posedge WCLK, negedge WADDR[3], 1.0);
   $setup(posedge WADDR[4], posedge WCLK, 1.0);
   $setup(negedge WADDR[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[4], 1.0);
   $hold(posedge WCLK, negedge WADDR[4], 1.0);
   $setup(posedge WADDR[5], posedge WCLK, 1.0);
   $setup(negedge WADDR[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[5], 1.0);
   $hold(posedge WCLK, negedge WADDR[5], 1.0);
   $setup(posedge WADDR[6], posedge WCLK, 1.0);
   $setup(negedge WADDR[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[6], 1.0);
   $hold(posedge WCLK, negedge WADDR[6], 1.0);
   $setup(posedge WADDR[7], posedge WCLK, 1.0);
   $setup(negedge WADDR[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[7], 1.0);
   $hold(posedge WCLK, negedge WADDR[7], 1.0);
   $setup(posedge WADDR[8], posedge WCLK, 1.0);
   $setup(negedge WADDR[8], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[8], 1.0);
   $hold(posedge WCLK, negedge WADDR[8], 1.0);
   $setup(posedge WADDR[9], posedge WCLK, 1.0);
   $setup(negedge WADDR[9], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[9], 1.0);
   $hold(posedge WCLK, negedge WADDR[9], 1.0);
   $setup(posedge WADDR[10], posedge WCLK, 1.0);
   $setup(negedge WADDR[10], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[10], 1.0);
   $hold(posedge WCLK, negedge WADDR[10], 1.0);
   $setup(posedge WADDR[11], posedge WCLK, 1.0);
   $setup(negedge WADDR[11], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[11], 1.0);
   $hold(posedge WCLK, negedge WADDR[11], 1.0);
   $setup(posedge WDATA[0], posedge WCLK, 1.0);
   $setup(negedge WDATA[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[0], 1.0);
   $hold(posedge WCLK, negedge WDATA[0], 1.0);
   $setup(posedge WDATA[1], posedge WCLK, 1.0);
   $setup(negedge WDATA[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[1], 1.0);
   $hold(posedge WCLK, negedge WDATA[1], 1.0);
   $setup(posedge WDATA[2], posedge WCLK, 1.0);
   $setup(negedge WDATA[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[2], 1.0);
   $hold(posedge WCLK, negedge WDATA[2], 1.0);
   $setup(posedge WDATA[3], posedge WCLK, 1.0);
   $setup(negedge WDATA[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[3], 1.0);
   $hold(posedge WCLK, negedge WDATA[3], 1.0);
   $setup(posedge WCLKE, posedge WCLK, 1.0);
   $setup(negedge WCLKE, posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WCLKE, 1.0);
   $hold(posedge WCLK, negedge WCLKE, 1.0);
   $setup(posedge WE, posedge WCLK, 1.0);
   $setup(negedge WE, posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WE, 1.0);
   $hold(posedge WCLK, negedge WE, 1.0);
   $setup(posedge RADDR[0], posedge RCLKN, 1.0);
   $setup(negedge RADDR[0], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[0], 1.0);
   $hold(posedge RCLKN, negedge RADDR[0], 1.0);
   $setup(posedge RADDR[1], posedge RCLKN, 1.0);
   $setup(negedge RADDR[1], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[1], 1.0);
   $hold(posedge RCLKN, negedge RADDR[1], 1.0);
   $setup(posedge RADDR[2], posedge RCLKN, 1.0);
   $setup(negedge RADDR[2], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[2], 1.0);
   $hold(posedge RCLKN, negedge RADDR[2], 1.0);
   $setup(posedge RADDR[3], posedge RCLKN, 1.0);
   $setup(negedge RADDR[3], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[3], 1.0);
   $hold(posedge RCLKN, negedge RADDR[3], 1.0);
   $setup(posedge RADDR[4], posedge RCLKN, 1.0);
   $setup(negedge RADDR[4], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[4], 1.0);
   $hold(posedge RCLKN, negedge RADDR[4], 1.0);
   $setup(posedge RADDR[5], posedge RCLKN, 1.0);
   $setup(negedge RADDR[5], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[5], 1.0);
   $hold(posedge RCLKN, negedge RADDR[5], 1.0);
   $setup(posedge RADDR[6], posedge RCLKN, 1.0);
   $setup(negedge RADDR[6], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[6], 1.0);
   $hold(posedge RCLKN, negedge RADDR[6], 1.0);
   $setup(posedge RADDR[7], posedge RCLKN, 1.0);
   $setup(negedge RADDR[7], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[7], 1.0);
   $hold(posedge RCLKN, negedge RADDR[7], 1.0);
   $setup(posedge RADDR[8], posedge RCLKN, 1.0);
   $setup(negedge RADDR[8], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[8], 1.0);
   $hold(posedge RCLKN, negedge RADDR[8], 1.0);
   $setup(posedge RADDR[9], posedge RCLKN, 1.0);
   $setup(negedge RADDR[9], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[9], 1.0);
   $hold(posedge RCLKN, negedge RADDR[9], 1.0);
   $setup(posedge RADDR[10], posedge RCLKN, 1.0);
   $setup(negedge RADDR[10], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[10], 1.0);
   $hold(posedge RCLKN, negedge RADDR[10], 1.0);
   $setup(posedge RADDR[11], posedge RCLKN, 1.0);
   $setup(negedge RADDR[11], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[11], 1.0);
   $hold(posedge RCLKN, negedge RADDR[11], 1.0);
   $setup(posedge RCLKE, posedge RCLKN, 1.0);
   $setup(negedge RCLKE, posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RCLKE, 1.0);
   $hold(posedge RCLKN, negedge RCLKE, 1.0);
   $setup(posedge RE, posedge RCLKN, 1.0);
   $setup(negedge RE, posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RE, 1.0);
   $hold(posedge RCLKN, negedge RE, 1.0);
endspecify
`endif
  
endmodule // SB_RAM4096x4NR 

//---------------------------------------
//	--- SB_RAM4096x4NW
//---------------------------------------
`timescale 1ps/1ps
module  SB_RAM4096x4NW ( RDATA, RCLK, RCLKE, RE, RADDR, WCLKN, WCLKE, WE, WADDR, WDATA ); 

output	[3:0]	RDATA;  
input         	RCLK;   
input           RCLKE; 
input           RE; 
input	[11:0]  RADDR; 
input           WCLKN; 
input           WCLKE; 
input           WE; 
input 	[11:0]  WADDR; 
input 	[3:0]	WDATA;

parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;


wire WCLK;
assign (weak0, weak1) RCLKE =1'b1 ;
assign (weak0, weak1) RE =1'b0 ;
assign (weak0, weak1) WCLKE =1'b1 ;
assign (weak0, weak1) WE =1'b0 ;
assign WCLK = ~WCLKN;

SB_RAM4096x4 sb_ram4096x4w_inst (
	.RDATA(RDATA),
	.RCLK(RCLK),
	.RCLKE(RCLKE),
	.RE(RE),
	.RADDR(RADDR),
	.WCLK(WCLK),
	.WCLKE(WCLKE),
	.WE(WE),
	.WADDR(WADDR),
	.WDATA(WDATA));

defparam sb_ram4096x4w_inst.INIT_0 = INIT_0;
defparam sb_ram4096x4w_inst.INIT_1 = INIT_1;
defparam sb_ram4096x4w_inst.INIT_2 = INIT_2;
defparam sb_ram4096x4w_inst.INIT_3 = INIT_3;
defparam sb_ram4096x4w_inst.INIT_4 = INIT_4;
defparam sb_ram4096x4w_inst.INIT_5 = INIT_5;
defparam sb_ram4096x4w_inst.INIT_6 = INIT_6;
defparam sb_ram4096x4w_inst.INIT_7 = INIT_7;
defparam sb_ram4096x4w_inst.INIT_8 = INIT_8;
defparam sb_ram4096x4w_inst.INIT_9 = INIT_9;
defparam sb_ram4096x4w_inst.INIT_A = INIT_A;
defparam sb_ram4096x4w_inst.INIT_B = INIT_B;
defparam sb_ram4096x4w_inst.INIT_C = INIT_C;
defparam sb_ram4096x4w_inst.INIT_D = INIT_D;
defparam sb_ram4096x4w_inst.INIT_E = INIT_E;
defparam sb_ram4096x4w_inst.INIT_F = INIT_F;

defparam sb_ram4096x4w_inst.INIT_10 = INIT_10;
defparam sb_ram4096x4w_inst.INIT_11 = INIT_11;
defparam sb_ram4096x4w_inst.INIT_12 = INIT_12;
defparam sb_ram4096x4w_inst.INIT_13 = INIT_13;
defparam sb_ram4096x4w_inst.INIT_14 = INIT_14;
defparam sb_ram4096x4w_inst.INIT_15 = INIT_15;
defparam sb_ram4096x4w_inst.INIT_16 = INIT_16;
defparam sb_ram4096x4w_inst.INIT_17 = INIT_17;
defparam sb_ram4096x4w_inst.INIT_18 = INIT_18;
defparam sb_ram4096x4w_inst.INIT_19 = INIT_19;
defparam sb_ram4096x4w_inst.INIT_1A = INIT_1A;
defparam sb_ram4096x4w_inst.INIT_1B = INIT_1B;
defparam sb_ram4096x4w_inst.INIT_1C = INIT_1C;
defparam sb_ram4096x4w_inst.INIT_1D = INIT_1D;
defparam sb_ram4096x4w_inst.INIT_1E = INIT_1E;
defparam sb_ram4096x4w_inst.INIT_1F = INIT_1F;

defparam sb_ram4096x4w_inst.INIT_20 = INIT_20;
defparam sb_ram4096x4w_inst.INIT_21 = INIT_21;
defparam sb_ram4096x4w_inst.INIT_22 = INIT_22;
defparam sb_ram4096x4w_inst.INIT_23 = INIT_23;
defparam sb_ram4096x4w_inst.INIT_24 = INIT_24;
defparam sb_ram4096x4w_inst.INIT_25 = INIT_25;
defparam sb_ram4096x4w_inst.INIT_26 = INIT_26;
defparam sb_ram4096x4w_inst.INIT_27 = INIT_27;
defparam sb_ram4096x4w_inst.INIT_28 = INIT_28;
defparam sb_ram4096x4w_inst.INIT_29 = INIT_29;
defparam sb_ram4096x4w_inst.INIT_2A = INIT_2A;
defparam sb_ram4096x4w_inst.INIT_2B = INIT_2B;
defparam sb_ram4096x4w_inst.INIT_2C = INIT_2C;
defparam sb_ram4096x4w_inst.INIT_2D = INIT_2D;
defparam sb_ram4096x4w_inst.INIT_2E = INIT_2E;
defparam sb_ram4096x4w_inst.INIT_2F = INIT_2F;

defparam sb_ram4096x4w_inst.INIT_30 = INIT_30;
defparam sb_ram4096x4w_inst.INIT_31 = INIT_31;
defparam sb_ram4096x4w_inst.INIT_32 = INIT_32;
defparam sb_ram4096x4w_inst.INIT_33 = INIT_33;
defparam sb_ram4096x4w_inst.INIT_34 = INIT_34;
defparam sb_ram4096x4w_inst.INIT_35 = INIT_35;
defparam sb_ram4096x4w_inst.INIT_36 = INIT_36;
defparam sb_ram4096x4w_inst.INIT_37 = INIT_37;
defparam sb_ram4096x4w_inst.INIT_38 = INIT_38;
defparam sb_ram4096x4w_inst.INIT_39 = INIT_39;
defparam sb_ram4096x4w_inst.INIT_3A = INIT_3A;
defparam sb_ram4096x4w_inst.INIT_3B = INIT_3B;
defparam sb_ram4096x4w_inst.INIT_3C = INIT_3C;
defparam sb_ram4096x4w_inst.INIT_3D = INIT_3D;
defparam sb_ram4096x4w_inst.INIT_3E = INIT_3E;
defparam sb_ram4096x4w_inst.INIT_3F = INIT_3F;


`ifdef TIMINGCHECK
specify
   (RCLK *> RDATA[0]) = (1.0, 1.0);
   (RCLK *> RDATA[1]) = (1.0, 1.0);
   (RCLK *> RDATA[2]) = (1.0, 1.0);
   (RCLK *> RDATA[3]) = (1.0, 1.0);
   $setup(posedge WADDR[0], posedge WCLKN, 1.0);
   $setup(negedge WADDR[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[0], 1.0);
   $hold(posedge WCLKN, negedge WADDR[0], 1.0);
   $setup(posedge WADDR[1], posedge WCLKN, 1.0);
   $setup(negedge WADDR[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[1], 1.0);
   $hold(posedge WCLKN, negedge WADDR[1], 1.0);
   $setup(posedge WADDR[2], posedge WCLKN, 1.0);
   $setup(negedge WADDR[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[2], 1.0);
   $hold(posedge WCLKN, negedge WADDR[2], 1.0);
   $setup(posedge WADDR[3], posedge WCLKN, 1.0);
   $setup(negedge WADDR[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[3], 1.0);
   $hold(posedge WCLKN, negedge WADDR[3], 1.0);
   $setup(posedge WADDR[4], posedge WCLKN, 1.0);
   $setup(negedge WADDR[4], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[4], 1.0);
   $hold(posedge WCLKN, negedge WADDR[4], 1.0);
   $setup(posedge WADDR[5], posedge WCLKN, 1.0);
   $setup(negedge WADDR[5], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[5], 1.0);
   $hold(posedge WCLKN, negedge WADDR[5], 1.0);
   $setup(posedge WADDR[6], posedge WCLKN, 1.0);
   $setup(negedge WADDR[6], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[6], 1.0);
   $hold(posedge WCLKN, negedge WADDR[6], 1.0);
   $setup(posedge WADDR[7], posedge WCLKN, 1.0);
   $setup(negedge WADDR[7], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[7], 1.0);
   $hold(posedge WCLKN, negedge WADDR[7], 1.0);
   $setup(posedge WADDR[8], posedge WCLKN, 1.0);
   $setup(negedge WADDR[8], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[8], 1.0);
   $hold(posedge WCLKN, negedge WADDR[8], 1.0);
   $setup(posedge WADDR[9], posedge WCLKN, 1.0);
   $setup(negedge WADDR[9], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[9], 1.0);
   $hold(posedge WCLKN, negedge WADDR[9], 1.0);
   $setup(posedge WADDR[10], posedge WCLKN, 1.0);
   $setup(negedge WADDR[10], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[10], 1.0);
   $hold(posedge WCLKN, negedge WADDR[10], 1.0);
   $setup(posedge WADDR[11], posedge WCLKN, 1.0);
   $setup(negedge WADDR[11], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[11], 1.0);
   $hold(posedge WCLKN, negedge WADDR[11], 1.0);
   $setup(posedge WDATA[0], posedge WCLKN, 1.0);
   $setup(negedge WDATA[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[0], 1.0);
   $hold(posedge WCLKN, negedge WDATA[0], 1.0);
   $setup(posedge WDATA[1], posedge WCLKN, 1.0);
   $setup(negedge WDATA[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[1], 1.0);
   $hold(posedge WCLKN, negedge WDATA[1], 1.0);
   $setup(posedge WDATA[2], posedge WCLKN, 1.0);
   $setup(negedge WDATA[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[2], 1.0);
   $hold(posedge WCLKN, negedge WDATA[2], 1.0);
   $setup(posedge WDATA[3], posedge WCLKN, 1.0);
   $setup(negedge WDATA[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[3], 1.0);
   $hold(posedge WCLKN, negedge WDATA[3], 1.0);
   $setup(posedge WCLKE, posedge WCLKN, 1.0);
   $setup(negedge WCLKE, posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WCLKE, 1.0);
   $hold(posedge WCLKN, negedge WCLKE, 1.0);
   $setup(posedge WE, posedge WCLKN, 1.0);
   $setup(negedge WE, posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WE, 1.0);
   $hold(posedge WCLKN, negedge WE, 1.0);
   $setup(posedge RADDR[0], posedge RCLK, 1.0);
   $setup(negedge RADDR[0], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[0], 1.0);
   $hold(posedge RCLK, negedge RADDR[0], 1.0);
   $setup(posedge RADDR[1], posedge RCLK, 1.0);
   $setup(negedge RADDR[1], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[1], 1.0);
   $hold(posedge RCLK, negedge RADDR[1], 1.0);
   $setup(posedge RADDR[2], posedge RCLK, 1.0);
   $setup(negedge RADDR[2], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[2], 1.0);
   $hold(posedge RCLK, negedge RADDR[2], 1.0);
   $setup(posedge RADDR[3], posedge RCLK, 1.0);
   $setup(negedge RADDR[3], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[3], 1.0);
   $hold(posedge RCLK, negedge RADDR[3], 1.0);
   $setup(posedge RADDR[4], posedge RCLK, 1.0);
   $setup(negedge RADDR[4], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[4], 1.0);
   $hold(posedge RCLK, negedge RADDR[4], 1.0);
   $setup(posedge RADDR[5], posedge RCLK, 1.0);
   $setup(negedge RADDR[5], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[5], 1.0);
   $hold(posedge RCLK, negedge RADDR[5], 1.0);
   $setup(posedge RADDR[6], posedge RCLK, 1.0);
   $setup(negedge RADDR[6], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[6], 1.0);
   $hold(posedge RCLK, negedge RADDR[6], 1.0);
   $setup(posedge RADDR[7], posedge RCLK, 1.0);
   $setup(negedge RADDR[7], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[7], 1.0);
   $hold(posedge RCLK, negedge RADDR[7], 1.0);
   $setup(posedge RADDR[8], posedge RCLK, 1.0);
   $setup(negedge RADDR[8], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[8], 1.0);
   $hold(posedge RCLK, negedge RADDR[8], 1.0);
   $setup(posedge RADDR[9], posedge RCLK, 1.0);
   $setup(negedge RADDR[9], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[9], 1.0);
   $hold(posedge RCLK, negedge RADDR[9], 1.0);
   $setup(posedge RADDR[10], posedge RCLK, 1.0);
   $setup(negedge RADDR[10], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[10], 1.0);
   $hold(posedge RCLK, negedge RADDR[10], 1.0);
   $setup(posedge RADDR[11], posedge RCLK, 1.0);
   $setup(negedge RADDR[11], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[11], 1.0);
   $hold(posedge RCLK, negedge RADDR[11], 1.0);
   $setup(posedge RCLKE, posedge RCLK, 1.0);
   $setup(negedge RCLKE, posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RCLKE, 1.0);
   $hold(posedge RCLK, negedge RCLKE, 1.0);
   $setup(posedge RE, posedge RCLK, 1.0);
   $setup(negedge RE, posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RE, 1.0);
   $hold(posedge RCLK, negedge RE, 1.0);
endspecify
`endif

endmodule  	// SB_RAM4096x4NW

//---------------------------------------
//	--- SB_RAM4096x4NRNW
//---------------------------------------
`timescale 1ps/1ps
module SB_RAM4096x4NRNW ( RDATA, RCLKN, RCLKE, RE, RADDR, WCLKN, WCLKE, WE, WADDR, WDATA ); 

output	[3:0]	RDATA;  
input         	RCLKN;   
input           RCLKE; 
input           RE; 
input	[11:0]  RADDR; 
input           WCLKN; 
input           WCLKE; 
input           WE; 
input 	[11:0]  WADDR; 
input 	[3:0]	WDATA;
  
parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;


wire RCLK, WCLK;
assign (weak0, weak1) RCLKE =1'b1 ;
assign (weak0, weak1) RE =1'b0 ;
assign (weak0, weak1) WCLKE =1'b1 ;
assign (weak0, weak1) WE =1'b0 ;
assign RCLK = ~RCLKN;
assign WCLK = ~WCLKN;

SB_RAM4096x4 sb_ram4096x4rw_inst (
	.RDATA(RDATA),
	.RCLK(RCLK),
	.RCLKE(RCLKE),
	.RE(RE),
	.RADDR(RADDR),
	.WCLK(WCLK),
	.WCLKE(WCLKE),
	.WE(WE),
	.WADDR(WADDR),
	.WDATA(WDATA));

defparam sb_ram4096x4rw_inst.INIT_0 = INIT_0;
defparam sb_ram4096x4rw_inst.INIT_1 = INIT_1;
defparam sb_ram4096x4rw_inst.INIT_2 = INIT_2;
defparam sb_ram4096x4rw_inst.INIT_3 = INIT_3;
defparam sb_ram4096x4rw_inst.INIT_4 = INIT_4;
defparam sb_ram4096x4rw_inst.INIT_5 = INIT_5;
defparam sb_ram4096x4rw_inst.INIT_6 = INIT_6;
defparam sb_ram4096x4rw_inst.INIT_7 = INIT_7;
defparam sb_ram4096x4rw_inst.INIT_8 = INIT_8;
defparam sb_ram4096x4rw_inst.INIT_9 = INIT_9;
defparam sb_ram4096x4rw_inst.INIT_A = INIT_A;
defparam sb_ram4096x4rw_inst.INIT_B = INIT_B;
defparam sb_ram4096x4rw_inst.INIT_C = INIT_C;
defparam sb_ram4096x4rw_inst.INIT_D = INIT_D;
defparam sb_ram4096x4rw_inst.INIT_E = INIT_E;
defparam sb_ram4096x4rw_inst.INIT_F = INIT_F;

defparam sb_ram4096x4rw_inst.INIT_10 = INIT_10;
defparam sb_ram4096x4rw_inst.INIT_11 = INIT_11;
defparam sb_ram4096x4rw_inst.INIT_12 = INIT_12;
defparam sb_ram4096x4rw_inst.INIT_13 = INIT_13;
defparam sb_ram4096x4rw_inst.INIT_14 = INIT_14;
defparam sb_ram4096x4rw_inst.INIT_15 = INIT_15;
defparam sb_ram4096x4rw_inst.INIT_16 = INIT_16;
defparam sb_ram4096x4rw_inst.INIT_17 = INIT_17;
defparam sb_ram4096x4rw_inst.INIT_18 = INIT_18;
defparam sb_ram4096x4rw_inst.INIT_19 = INIT_19;
defparam sb_ram4096x4rw_inst.INIT_1A = INIT_1A;
defparam sb_ram4096x4rw_inst.INIT_1B = INIT_1B;
defparam sb_ram4096x4rw_inst.INIT_1C = INIT_1C;
defparam sb_ram4096x4rw_inst.INIT_1D = INIT_1D;
defparam sb_ram4096x4rw_inst.INIT_1E = INIT_1E;
defparam sb_ram4096x4rw_inst.INIT_1F = INIT_1F;

defparam sb_ram4096x4rw_inst.INIT_20 = INIT_20;
defparam sb_ram4096x4rw_inst.INIT_21 = INIT_21;
defparam sb_ram4096x4rw_inst.INIT_22 = INIT_22;
defparam sb_ram4096x4rw_inst.INIT_23 = INIT_23;
defparam sb_ram4096x4rw_inst.INIT_24 = INIT_24;
defparam sb_ram4096x4rw_inst.INIT_25 = INIT_25;
defparam sb_ram4096x4rw_inst.INIT_26 = INIT_26;
defparam sb_ram4096x4rw_inst.INIT_27 = INIT_27;
defparam sb_ram4096x4rw_inst.INIT_28 = INIT_28;
defparam sb_ram4096x4rw_inst.INIT_29 = INIT_29;
defparam sb_ram4096x4rw_inst.INIT_2A = INIT_2A;
defparam sb_ram4096x4rw_inst.INIT_2B = INIT_2B;
defparam sb_ram4096x4rw_inst.INIT_2C = INIT_2C;
defparam sb_ram4096x4rw_inst.INIT_2D = INIT_2D;
defparam sb_ram4096x4rw_inst.INIT_2E = INIT_2E;
defparam sb_ram4096x4rw_inst.INIT_2F = INIT_2F;

defparam sb_ram4096x4rw_inst.INIT_30 = INIT_30;
defparam sb_ram4096x4rw_inst.INIT_31 = INIT_31;
defparam sb_ram4096x4rw_inst.INIT_32 = INIT_32;
defparam sb_ram4096x4rw_inst.INIT_33 = INIT_33;
defparam sb_ram4096x4rw_inst.INIT_34 = INIT_34;
defparam sb_ram4096x4rw_inst.INIT_35 = INIT_35;
defparam sb_ram4096x4rw_inst.INIT_36 = INIT_36;
defparam sb_ram4096x4rw_inst.INIT_37 = INIT_37;
defparam sb_ram4096x4rw_inst.INIT_38 = INIT_38;
defparam sb_ram4096x4rw_inst.INIT_39 = INIT_39;
defparam sb_ram4096x4rw_inst.INIT_3A = INIT_3A;
defparam sb_ram4096x4rw_inst.INIT_3B = INIT_3B;
defparam sb_ram4096x4rw_inst.INIT_3C = INIT_3C;
defparam sb_ram4096x4rw_inst.INIT_3D = INIT_3D;
defparam sb_ram4096x4rw_inst.INIT_3E = INIT_3E;
defparam sb_ram4096x4rw_inst.INIT_3F = INIT_3F;


`ifdef TIMINGCHECK
specify
   (RCLKN *> RDATA[0]) = (1.0, 1.0);
   (RCLKN *> RDATA[1]) = (1.0, 1.0);
   (RCLKN *> RDATA[2]) = (1.0, 1.0);
   (RCLKN *> RDATA[3]) = (1.0, 1.0);
   $setup(posedge WADDR[0], posedge WCLKN, 1.0);
   $setup(negedge WADDR[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[0], 1.0);
   $hold(posedge WCLKN, negedge WADDR[0], 1.0);
   $setup(posedge WADDR[1], posedge WCLKN, 1.0);
   $setup(negedge WADDR[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[1], 1.0);
   $hold(posedge WCLKN, negedge WADDR[1], 1.0);
   $setup(posedge WADDR[2], posedge WCLKN, 1.0);
   $setup(negedge WADDR[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[2], 1.0);
   $hold(posedge WCLKN, negedge WADDR[2], 1.0);
   $setup(posedge WADDR[3], posedge WCLKN, 1.0);
   $setup(negedge WADDR[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[3], 1.0);
   $hold(posedge WCLKN, negedge WADDR[3], 1.0);
   $setup(posedge WADDR[4], posedge WCLKN, 1.0);
   $setup(negedge WADDR[4], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[4], 1.0);
   $hold(posedge WCLKN, negedge WADDR[4], 1.0);
   $setup(posedge WADDR[5], posedge WCLKN, 1.0);
   $setup(negedge WADDR[5], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[5], 1.0);
   $hold(posedge WCLKN, negedge WADDR[5], 1.0);
   $setup(posedge WADDR[6], posedge WCLKN, 1.0);
   $setup(negedge WADDR[6], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[6], 1.0);
   $hold(posedge WCLKN, negedge WADDR[6], 1.0);
   $setup(posedge WADDR[7], posedge WCLKN, 1.0);
   $setup(negedge WADDR[7], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[7], 1.0);
   $hold(posedge WCLKN, negedge WADDR[7], 1.0);
   $setup(posedge WADDR[8], posedge WCLKN, 1.0);
   $setup(negedge WADDR[8], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[8], 1.0);
   $hold(posedge WCLKN, negedge WADDR[8], 1.0);
   $setup(posedge WADDR[9], posedge WCLKN, 1.0);
   $setup(negedge WADDR[9], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[9], 1.0);
   $hold(posedge WCLKN, negedge WADDR[9], 1.0);
   $setup(posedge WADDR[10], posedge WCLKN, 1.0);
   $setup(negedge WADDR[10], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[10], 1.0);
   $hold(posedge WCLKN, negedge WADDR[10], 1.0);
   $setup(posedge WADDR[11], posedge WCLKN, 1.0);
   $setup(negedge WADDR[11], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[11], 1.0);
   $hold(posedge WCLKN, negedge WADDR[11], 1.0);
   $setup(posedge WDATA[0], posedge WCLKN, 1.0);
   $setup(negedge WDATA[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[0], 1.0);
   $hold(posedge WCLKN, negedge WDATA[0], 1.0);
   $setup(posedge WDATA[1], posedge WCLKN, 1.0);
   $setup(negedge WDATA[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[1], 1.0);
   $hold(posedge WCLKN, negedge WDATA[1], 1.0);
   $setup(posedge WDATA[2], posedge WCLKN, 1.0);
   $setup(negedge WDATA[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[2], 1.0);
   $hold(posedge WCLKN, negedge WDATA[2], 1.0);
   $setup(posedge WDATA[3], posedge WCLKN, 1.0);
   $setup(negedge WDATA[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[3], 1.0);
   $hold(posedge WCLKN, negedge WDATA[3], 1.0);
   $setup(posedge WCLKE, posedge WCLKN, 1.0);
   $setup(negedge WCLKE, posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WCLKE, 1.0);
   $hold(posedge WCLKN, negedge WCLKE, 1.0);
   $setup(posedge WE, posedge WCLKN, 1.0);
   $setup(negedge WE, posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WE, 1.0);
   $hold(posedge WCLKN, negedge WE, 1.0);
   $setup(posedge RADDR[0], posedge RCLKN, 1.0);
   $setup(negedge RADDR[0], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[0], 1.0);
   $hold(posedge RCLKN, negedge RADDR[0], 1.0);
   $setup(posedge RADDR[1], posedge RCLKN, 1.0);
   $setup(negedge RADDR[1], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[1], 1.0);
   $hold(posedge RCLKN, negedge RADDR[1], 1.0);
   $setup(posedge RADDR[2], posedge RCLKN, 1.0);
   $setup(negedge RADDR[2], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[2], 1.0);
   $hold(posedge RCLKN, negedge RADDR[2], 1.0);
   $setup(posedge RADDR[3], posedge RCLKN, 1.0);
   $setup(negedge RADDR[3], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[3], 1.0);
   $hold(posedge RCLKN, negedge RADDR[3], 1.0);
   $setup(posedge RADDR[4], posedge RCLKN, 1.0);
   $setup(negedge RADDR[4], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[4], 1.0);
   $hold(posedge RCLKN, negedge RADDR[4], 1.0);
   $setup(posedge RADDR[5], posedge RCLKN, 1.0);
   $setup(negedge RADDR[5], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[5], 1.0);
   $hold(posedge RCLKN, negedge RADDR[5], 1.0);
   $setup(posedge RADDR[6], posedge RCLKN, 1.0);
   $setup(negedge RADDR[6], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[6], 1.0);
   $hold(posedge RCLKN, negedge RADDR[6], 1.0);
   $setup(posedge RADDR[7], posedge RCLKN, 1.0);
   $setup(negedge RADDR[7], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[7], 1.0);
   $hold(posedge RCLKN, negedge RADDR[7], 1.0);
   $setup(posedge RADDR[8], posedge RCLKN, 1.0);
   $setup(negedge RADDR[8], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[8], 1.0);
   $hold(posedge RCLKN, negedge RADDR[8], 1.0);
   $setup(posedge RADDR[9], posedge RCLKN, 1.0);
   $setup(negedge RADDR[9], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[9], 1.0);
   $hold(posedge RCLKN, negedge RADDR[9], 1.0);
   $setup(posedge RADDR[10], posedge RCLKN, 1.0);
   $setup(negedge RADDR[10], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[10], 1.0);
   $hold(posedge RCLKN, negedge RADDR[10], 1.0);
   $setup(posedge RADDR[11], posedge RCLKN, 1.0);
   $setup(negedge RADDR[11], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[11], 1.0);
   $hold(posedge RCLKN, negedge RADDR[11], 1.0);
   $setup(posedge RCLKE, posedge RCLKN, 1.0);
   $setup(negedge RCLKE, posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RCLKE, 1.0);
   $hold(posedge RCLKN, negedge RCLKE, 1.0);
   $setup(posedge RE, posedge RCLKN, 1.0);
   $setup(negedge RE, posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RE, 1.0);
   $hold(posedge RCLKN, negedge RE, 1.0);
endspecify
`endif

endmodule 	// SB_RAM4096x4NRNW 

//---------------------------------------
//	--- SB_RAM8192x2
//---------------------------------------
`timescale 1ps/1ps
module SB_RAM8192x2  ( RDATA, RCLK, RCLKE, RE, RADDR, WCLK, WCLKE, WE, WADDR, WDATA ); 

output	[1:0]	RDATA;  
input         	RCLK;   
input           RCLKE; 
input           RE; 
input	[12:0]  RADDR; 
input           WCLK; 
input           WCLKE; 
input           WE; 
input 	[12:0]  WADDR; 
input 	[1:0]	WDATA; 
  
parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

// local Parameters
localparam			CLOCK_PERIOD = 200;	//
localparam 			DELAY	= (CLOCK_PERIOD/10);		// Clock-to-output delay. Zero
							// time delays can be confusing
							// and sometimes cause problems.
localparam 			BUS_WIDTH = 2;		// Width of RAM (number of bits)

localparam 			ADDRESS_BUS_SIZE = 13;	// Number of bits required to
							// represent the RAM address

localparam   ADDRESSABLE_SPACE  = 2**ADDRESS_BUS_SIZE;	// Decimal address range [2^Size:0]


// SIGNAL DECLARATIONS
wire			   	WCLK_g, RCLK_g;
reg 				WCLKE_sync, RCLKE_sync; 
assign (weak0, weak1) RCLKE =1'b1 ;
assign (weak0, weak1) RE =1'b0 ;
assign (weak0, weak1) WCLKE =1'b1 ;
assign (weak0, weak1) WE =1'b0 ;
reg	Memory	[BUS_WIDTH*ADDRESSABLE_SPACE-1:0];
// 
event Read_e, Write_e;

//////////////////// Collision detect begins here ///////////////////////////////
localparam 	TRUE = 1'b1;
localparam	FALSE = 1'b0;
reg 		Time_Collision_Detected = 1'b0;
wire		Address_Collision_Detected;

event Collision_e;

time COLLISION_TIME_WINDOW = (CLOCK_PERIOD/8); // This is an arbitray value, but is better than using an absolute 
						    // value, because the actual time window depends on the actual silicon 
						    // implementation. Thus the test is indicative of an Error and not
						    // guaranteed to be an error. Even so this is usefull.
time time_WCLK_RCLK, time_WCLK, time_RCLK;


//function reg Check_Timed_Window_Violation;
function	Check_Timed_Window_Violation;	
input T1, T2, Minimum_Time_Window;
time T1, T2;
time Minimum_Time_Window;
time Difference;	
	begin
		Difference = (T1 - T2);
		if (Difference < 0) Difference = -Difference;
		Check_Timed_Window_Violation = (Difference < Minimum_Time_Window);
	end
endfunction


initial begin
       time_WCLK = CLOCK_PERIOD;	// Arbitrary initialisation value, ensure no window collison error on first clock edge.
       time_RCLK = (CLOCK_PERIOD*8);	// Arbitrary initialisation difference value, ensure no collision error on first clock edge.					
end

integer	i,j;


initial	//	initialize ram_16k (8192 x 2) by init parameters, section by section
begin
	for	(i=0; i<=(256/BUS_WIDTH)-1; i=i+1)       
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)    
		begin 

			Memory[BUS_WIDTH*i+j]		=	INIT_0[BUS_WIDTH*i+j];
			Memory[256*1+BUS_WIDTH*i+j]	=	INIT_1[BUS_WIDTH*i+j];
			Memory[256*2+BUS_WIDTH*i+j]	=	INIT_2[BUS_WIDTH*i+j];
			Memory[256*3+BUS_WIDTH*i+j]	=	INIT_3[BUS_WIDTH*i+j];
			Memory[256*4+BUS_WIDTH*i+j]	=	INIT_4[BUS_WIDTH*i+j];
			Memory[256*5+BUS_WIDTH*i+j]	=	INIT_5[BUS_WIDTH*i+j];
			Memory[256*6+BUS_WIDTH*i+j]	=	INIT_6[BUS_WIDTH*i+j];
			Memory[256*7+BUS_WIDTH*i+j]	=	INIT_7[BUS_WIDTH*i+j];
			Memory[256*8+BUS_WIDTH*i+j]	=	INIT_8[BUS_WIDTH*i+j];
			Memory[256*9+BUS_WIDTH*i+j]	=	INIT_9[BUS_WIDTH*i+j];
			Memory[256*10+BUS_WIDTH*i+j]	=	INIT_A[BUS_WIDTH*i+j];
			Memory[256*11+BUS_WIDTH*i+j]	=	INIT_B[BUS_WIDTH*i+j];
			Memory[256*12+BUS_WIDTH*i+j]	=	INIT_C[BUS_WIDTH*i+j];
			Memory[256*13+BUS_WIDTH*i+j]	=	INIT_D[BUS_WIDTH*i+j];
			Memory[256*14+BUS_WIDTH*i+j]	=	INIT_E[BUS_WIDTH*i+j];
			Memory[256*15+BUS_WIDTH*i+j]	=	INIT_F[BUS_WIDTH*i+j];

			Memory[256*16+BUS_WIDTH*i+j]	=	INIT_10[BUS_WIDTH*i+j];
			Memory[256*17+BUS_WIDTH*i+j]	=	INIT_11[BUS_WIDTH*i+j];
			Memory[256*18+BUS_WIDTH*i+j]	=	INIT_12[BUS_WIDTH*i+j];
			Memory[256*19+BUS_WIDTH*i+j]	=	INIT_13[BUS_WIDTH*i+j];
			Memory[256*20+BUS_WIDTH*i+j]	=	INIT_14[BUS_WIDTH*i+j];
			Memory[256*21+BUS_WIDTH*i+j]	=	INIT_15[BUS_WIDTH*i+j];
			Memory[256*22+BUS_WIDTH*i+j]	=	INIT_16[BUS_WIDTH*i+j];
			Memory[256*23+BUS_WIDTH*i+j]	=	INIT_17[BUS_WIDTH*i+j];
			Memory[256*24+BUS_WIDTH*i+j]	=	INIT_18[BUS_WIDTH*i+j];
			Memory[256*25+BUS_WIDTH*i+j]	=	INIT_19[BUS_WIDTH*i+j];
			Memory[256*26+BUS_WIDTH*i+j]	=	INIT_1A[BUS_WIDTH*i+j];
			Memory[256*27+BUS_WIDTH*i+j]	=	INIT_1B[BUS_WIDTH*i+j];
			Memory[256*28+BUS_WIDTH*i+j]	=	INIT_1C[BUS_WIDTH*i+j];
			Memory[256*29+BUS_WIDTH*i+j]	=	INIT_1D[BUS_WIDTH*i+j];
			Memory[256*30+BUS_WIDTH*i+j]	=	INIT_1E[BUS_WIDTH*i+j];
			Memory[256*31+BUS_WIDTH*i+j]	=	INIT_1F[BUS_WIDTH*i+j];

			Memory[256*32+BUS_WIDTH*i+j]	=	INIT_20[BUS_WIDTH*i+j];
			Memory[256*33+BUS_WIDTH*i+j]	=	INIT_21[BUS_WIDTH*i+j];
			Memory[256*34+BUS_WIDTH*i+j]	=	INIT_22[BUS_WIDTH*i+j];
			Memory[256*35+BUS_WIDTH*i+j]	=	INIT_23[BUS_WIDTH*i+j];
			Memory[256*36+BUS_WIDTH*i+j]	=	INIT_24[BUS_WIDTH*i+j];
			Memory[256*37+BUS_WIDTH*i+j]	=	INIT_25[BUS_WIDTH*i+j];
			Memory[256*38+BUS_WIDTH*i+j]	=	INIT_26[BUS_WIDTH*i+j];
			Memory[256*39+BUS_WIDTH*i+j]	=	INIT_27[BUS_WIDTH*i+j];
			Memory[256*40+BUS_WIDTH*i+j]	=	INIT_28[BUS_WIDTH*i+j];
			Memory[256*41+BUS_WIDTH*i+j]	=	INIT_29[BUS_WIDTH*i+j];
			Memory[256*42+BUS_WIDTH*i+j]	=	INIT_2A[BUS_WIDTH*i+j];
			Memory[256*43+BUS_WIDTH*i+j]	=	INIT_2B[BUS_WIDTH*i+j];
			Memory[256*44+BUS_WIDTH*i+j]	=	INIT_2C[BUS_WIDTH*i+j];
			Memory[256*45+BUS_WIDTH*i+j]	=	INIT_2D[BUS_WIDTH*i+j];
			Memory[256*46+BUS_WIDTH*i+j]	=	INIT_2E[BUS_WIDTH*i+j];
			Memory[256*47+BUS_WIDTH*i+j]	=	INIT_2F[BUS_WIDTH*i+j];

			Memory[256*48+BUS_WIDTH*i+j]	=	INIT_30[BUS_WIDTH*i+j];
			Memory[256*49+BUS_WIDTH*i+j]	=	INIT_31[BUS_WIDTH*i+j];
			Memory[256*50+BUS_WIDTH*i+j]	=	INIT_32[BUS_WIDTH*i+j];
			Memory[256*51+BUS_WIDTH*i+j]	=	INIT_33[BUS_WIDTH*i+j];
			Memory[256*52+BUS_WIDTH*i+j]	=	INIT_34[BUS_WIDTH*i+j];
			Memory[256*53+BUS_WIDTH*i+j]	=	INIT_35[BUS_WIDTH*i+j];
			Memory[256*54+BUS_WIDTH*i+j]	=	INIT_36[BUS_WIDTH*i+j];
			Memory[256*55+BUS_WIDTH*i+j]	=	INIT_37[BUS_WIDTH*i+j];
			Memory[256*56+BUS_WIDTH*i+j]	=	INIT_38[BUS_WIDTH*i+j];
			Memory[256*57+BUS_WIDTH*i+j]	=	INIT_39[BUS_WIDTH*i+j];
			Memory[256*58+BUS_WIDTH*i+j]	=	INIT_3A[BUS_WIDTH*i+j];
			Memory[256*59+BUS_WIDTH*i+j]	=	INIT_3B[BUS_WIDTH*i+j];
			Memory[256*60+BUS_WIDTH*i+j]	=	INIT_3C[BUS_WIDTH*i+j];
			Memory[256*61+BUS_WIDTH*i+j]	=	INIT_3D[BUS_WIDTH*i+j];
			Memory[256*62+BUS_WIDTH*i+j]	=	INIT_3E[BUS_WIDTH*i+j];
			Memory[256*63+BUS_WIDTH*i+j]	=	INIT_3F[BUS_WIDTH*i+j];

		end 
	end

end

assign Address_Collision_Detected = ((RE & WE & WCLKE & RCLKE)&(WADDR == RADDR)); 

always @(WCLK or WCLKE) 
begin 
	if(~WCLK)
	WCLKE_sync = WCLKE;   	
end 

always @(RCLK or RCLKE) 
begin 
	if (~RCLK)
	RCLKE_sync = RCLKE; 	
end 

assign WCLK_g = WCLK & WCLKE_sync;
assign RCLK_g = RCLK & RCLKE_sync;


always @(posedge WCLK_g) begin
	time_WCLK = $time;
end

always @(posedge RCLK_g) begin
    	time_RCLK = $time;
end
integer	SB_RAM8192x2_RDATA_log_file;					//.....................
initial	SB_RAM8192x2_RDATA_log_file=("SB_RAM8192x2_RDATA_log_file.txt");	//.....................
always @(posedge WCLK_g) begin

	Time_Collision_Detected = Check_Timed_Window_Violation(time_WCLK,time_RCLK,COLLISION_TIME_WINDOW);
        if (Time_Collision_Detected & Address_Collision_Detected)begin
        	$display("Warning: Write-Read collision detected, Data read value is XXXX\n");
 		$display("WCLK Time: %.3f   RCLK Time:%.3f  ",time_WCLK, time_RCLK,"WADDR: %d   RADDR:%d\n",WADDR, RADDR); 
 		$fdisplay(SB_RAM8192x2_RDATA_log_file,"Warning: Write-Read collision detected, Data read value is XXXX\n");
		$fdisplay(SB_RAM8192x2_RDATA_log_file,"WCLK Time: %.3f   RCLK Time:%.3f  ",time_WCLK, time_RCLK, "WADDR: %d   RADDR:%d\n",WADDR, RADDR); 	
 		-> Collision_e;
	end
end

//	code modify for universal verilog compiler

always @ (posedge WCLK_g)
begin
	if	(WE)
	begin
		-> Write_e;
		for	(i=0;i<=BUS_WIDTH-1; i=i+1)
		begin
				Memory[WADDR*BUS_WIDTH+i]	<=	WDATA[i];
		end
	end
end

reg	[BUS_WIDTH-1:0]	RDATA = 0;

// Look at the rising edge of the clock

always @ (posedge RCLK_g)
begin
	if	(RE)
	begin
		-> Read_e;
		if	(Time_Collision_Detected & Address_Collision_Detected) 
			RDATA <= {BUS_WIDTH{1'hX}};
		else
			for	(i=0;i<=BUS_WIDTH-1;i=i+1)
				RDATA[i]	<= Memory[RADDR*BUS_WIDTH+i];
	end
end

`ifdef TIMINGCHECK
specify
   (RCLK *> RDATA[0]) = (1.0, 1.0);
   (RCLK *> RDATA[1]) = (1.0, 1.0);
   $setup(posedge WADDR[0], posedge WCLK, 1.0);
   $setup(negedge WADDR[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[0], 1.0);
   $hold(posedge WCLK, negedge WADDR[0], 1.0);
   $setup(posedge WADDR[1], posedge WCLK, 1.0);
   $setup(negedge WADDR[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[1], 1.0);
   $hold(posedge WCLK, negedge WADDR[1], 1.0);
   $setup(posedge WADDR[2], posedge WCLK, 1.0);
   $setup(negedge WADDR[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[2], 1.0);
   $hold(posedge WCLK, negedge WADDR[2], 1.0);
   $setup(posedge WADDR[3], posedge WCLK, 1.0);
   $setup(negedge WADDR[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[3], 1.0);
   $hold(posedge WCLK, negedge WADDR[3], 1.0);
   $setup(posedge WADDR[4], posedge WCLK, 1.0);
   $setup(negedge WADDR[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[4], 1.0);
   $hold(posedge WCLK, negedge WADDR[4], 1.0);
   $setup(posedge WADDR[5], posedge WCLK, 1.0);
   $setup(negedge WADDR[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[5], 1.0);
   $hold(posedge WCLK, negedge WADDR[5], 1.0);
   $setup(posedge WADDR[6], posedge WCLK, 1.0);
   $setup(negedge WADDR[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[6], 1.0);
   $hold(posedge WCLK, negedge WADDR[6], 1.0);
   $setup(posedge WADDR[7], posedge WCLK, 1.0);
   $setup(negedge WADDR[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[7], 1.0);
   $hold(posedge WCLK, negedge WADDR[7], 1.0);
   $setup(posedge WADDR[8], posedge WCLK, 1.0);
   $setup(negedge WADDR[8], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[8], 1.0);
   $hold(posedge WCLK, negedge WADDR[8], 1.0);
   $setup(posedge WADDR[9], posedge WCLK, 1.0);
   $setup(negedge WADDR[9], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[9], 1.0);
   $hold(posedge WCLK, negedge WADDR[9], 1.0);
   $setup(posedge WADDR[10], posedge WCLK, 1.0);
   $setup(negedge WADDR[10], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[10], 1.0);
   $hold(posedge WCLK, negedge WADDR[10], 1.0);
   $setup(posedge WADDR[11], posedge WCLK, 1.0);
   $setup(negedge WADDR[11], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[11], 1.0);
   $hold(posedge WCLK, negedge WADDR[11], 1.0);
   $setup(posedge WADDR[12], posedge WCLK, 1.0);
   $setup(negedge WADDR[12], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[12], 1.0);
   $hold(posedge WCLK, negedge WADDR[12], 1.0);
   $setup(posedge WDATA[0], posedge WCLK, 1.0);
   $setup(negedge WDATA[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[0], 1.0);
   $hold(posedge WCLK, negedge WDATA[0], 1.0);
   $setup(posedge WDATA[1], posedge WCLK, 1.0);
   $setup(negedge WDATA[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[1], 1.0);
   $hold(posedge WCLK, negedge WDATA[1], 1.0);
   $setup(posedge WCLKE, posedge WCLK, 1.0);
   $setup(negedge WCLKE, posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WCLKE, 1.0);
   $hold(posedge WCLK, negedge WCLKE, 1.0);
   $setup(posedge WE, posedge WCLK, 1.0);
   $setup(negedge WE, posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WE, 1.0);
   $hold(posedge WCLK, negedge WE, 1.0);
   $setup(posedge RADDR[0], posedge RCLK, 1.0);
   $setup(negedge RADDR[0], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[0], 1.0);
   $hold(posedge RCLK, negedge RADDR[0], 1.0);
   $setup(posedge RADDR[1], posedge RCLK, 1.0);
   $setup(negedge RADDR[1], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[1], 1.0);
   $hold(posedge RCLK, negedge RADDR[1], 1.0);
   $setup(posedge RADDR[2], posedge RCLK, 1.0);
   $setup(negedge RADDR[2], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[2], 1.0);
   $hold(posedge RCLK, negedge RADDR[2], 1.0);
   $setup(posedge RADDR[3], posedge RCLK, 1.0);
   $setup(negedge RADDR[3], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[3], 1.0);
   $hold(posedge RCLK, negedge RADDR[3], 1.0);
   $setup(posedge RADDR[4], posedge RCLK, 1.0);
   $setup(negedge RADDR[4], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[4], 1.0);
   $hold(posedge RCLK, negedge RADDR[4], 1.0);
   $setup(posedge RADDR[5], posedge RCLK, 1.0);
   $setup(negedge RADDR[5], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[5], 1.0);
   $hold(posedge RCLK, negedge RADDR[5], 1.0);
   $setup(posedge RADDR[6], posedge RCLK, 1.0);
   $setup(negedge RADDR[6], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[6], 1.0);
   $hold(posedge RCLK, negedge RADDR[6], 1.0);
   $setup(posedge RADDR[7], posedge RCLK, 1.0);
   $setup(negedge RADDR[7], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[7], 1.0);
   $hold(posedge RCLK, negedge RADDR[7], 1.0);
   $setup(posedge RADDR[8], posedge RCLK, 1.0);
   $setup(negedge RADDR[8], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[8], 1.0);
   $hold(posedge RCLK, negedge RADDR[8], 1.0);
   $setup(posedge RADDR[9], posedge RCLK, 1.0);
   $setup(negedge RADDR[9], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[9], 1.0);
   $hold(posedge RCLK, negedge RADDR[9], 1.0);
   $setup(posedge RADDR[10], posedge RCLK, 1.0);
   $setup(negedge RADDR[10], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[10], 1.0);
   $hold(posedge RCLK, negedge RADDR[10], 1.0);
   $setup(posedge RADDR[11], posedge RCLK, 1.0);
   $setup(negedge RADDR[11], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[11], 1.0);
   $hold(posedge RCLK, negedge RADDR[11], 1.0);
   $setup(posedge RADDR[12], posedge RCLK, 1.0);
   $setup(negedge RADDR[12], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[12], 1.0);
   $hold(posedge RCLK, negedge RADDR[12], 1.0);
   $setup(posedge RCLKE, posedge RCLK, 1.0);
   $setup(negedge RCLKE, posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RCLKE, 1.0);
   $hold(posedge RCLK, negedge RCLKE, 1.0);
   $setup(posedge RE, posedge RCLK, 1.0);
   $setup(negedge RE, posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RE, 1.0);
   $hold(posedge RCLK, negedge RE, 1.0);
endspecify
`endif

endmodule // SB_RAM8192x2

//---------------------------------------
//	--- SB_RAM8192x2NR
//---------------------------------------
`timescale 1ps/1ps
module SB_RAM8192x2NR ( RDATA, RCLKN, RCLKE, RE, RADDR, WCLK, WCLKE, WE, WADDR, WDATA ); 

output	[1:0]	RDATA;  
input         	RCLKN;   
input           RCLKE; 
input           RE; 
input	[12:0]  RADDR; 
input           WCLK; 
input           WCLKE; 
input           WE; 
input 	[12:0]  WADDR; 
input 	[1:0]	WDATA;  

parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

wire RCLK;
assign (weak0, weak1) RCLKE =1'b1 ;
assign (weak0, weak1) RE =1'b0 ;
assign (weak0, weak1) WCLKE =1'b1 ;
assign (weak0, weak1) WE =1'b0 ;
assign RCLK = ~RCLKN;

SB_RAM8192x2 sb_ram8192x2r_inst (
	.RDATA(RDATA),
	.RCLK(RCLK),
	.RCLKE(RCLKE),
	.RE(RE),
	.RADDR(RADDR),
	.WCLK(WCLK),
	.WCLKE(WCLKE),
	.WE(WE),
	.WADDR(WADDR),
	.WDATA(WDATA));

defparam sb_ram8192x2r_inst.INIT_0 = INIT_0;
defparam sb_ram8192x2r_inst.INIT_1 = INIT_1;
defparam sb_ram8192x2r_inst.INIT_2 = INIT_2;
defparam sb_ram8192x2r_inst.INIT_3 = INIT_3;
defparam sb_ram8192x2r_inst.INIT_4 = INIT_4;
defparam sb_ram8192x2r_inst.INIT_5 = INIT_5;
defparam sb_ram8192x2r_inst.INIT_6 = INIT_6;
defparam sb_ram8192x2r_inst.INIT_7 = INIT_7;
defparam sb_ram8192x2r_inst.INIT_8 = INIT_8;
defparam sb_ram8192x2r_inst.INIT_9 = INIT_9;
defparam sb_ram8192x2r_inst.INIT_A = INIT_A;
defparam sb_ram8192x2r_inst.INIT_B = INIT_B;
defparam sb_ram8192x2r_inst.INIT_C = INIT_C;
defparam sb_ram8192x2r_inst.INIT_D = INIT_D;
defparam sb_ram8192x2r_inst.INIT_E = INIT_E;
defparam sb_ram8192x2r_inst.INIT_F = INIT_F;

defparam sb_ram8192x2r_inst.INIT_10 = INIT_10;
defparam sb_ram8192x2r_inst.INIT_11 = INIT_11;
defparam sb_ram8192x2r_inst.INIT_12 = INIT_12;
defparam sb_ram8192x2r_inst.INIT_13 = INIT_13;
defparam sb_ram8192x2r_inst.INIT_14 = INIT_14;
defparam sb_ram8192x2r_inst.INIT_15 = INIT_15;
defparam sb_ram8192x2r_inst.INIT_16 = INIT_16;
defparam sb_ram8192x2r_inst.INIT_17 = INIT_17;
defparam sb_ram8192x2r_inst.INIT_18 = INIT_18;
defparam sb_ram8192x2r_inst.INIT_19 = INIT_19;
defparam sb_ram8192x2r_inst.INIT_1A = INIT_1A;
defparam sb_ram8192x2r_inst.INIT_1B = INIT_1B;
defparam sb_ram8192x2r_inst.INIT_1C = INIT_1C;
defparam sb_ram8192x2r_inst.INIT_1D = INIT_1D;
defparam sb_ram8192x2r_inst.INIT_1E = INIT_1E;
defparam sb_ram8192x2r_inst.INIT_1F = INIT_1F;

defparam sb_ram8192x2r_inst.INIT_20 = INIT_20;
defparam sb_ram8192x2r_inst.INIT_21 = INIT_21;
defparam sb_ram8192x2r_inst.INIT_22 = INIT_22;
defparam sb_ram8192x2r_inst.INIT_23 = INIT_23;
defparam sb_ram8192x2r_inst.INIT_24 = INIT_24;
defparam sb_ram8192x2r_inst.INIT_25 = INIT_25;
defparam sb_ram8192x2r_inst.INIT_26 = INIT_26;
defparam sb_ram8192x2r_inst.INIT_27 = INIT_27;
defparam sb_ram8192x2r_inst.INIT_28 = INIT_28;
defparam sb_ram8192x2r_inst.INIT_29 = INIT_29;
defparam sb_ram8192x2r_inst.INIT_2A = INIT_2A;
defparam sb_ram8192x2r_inst.INIT_2B = INIT_2B;
defparam sb_ram8192x2r_inst.INIT_2C = INIT_2C;
defparam sb_ram8192x2r_inst.INIT_2D = INIT_2D;
defparam sb_ram8192x2r_inst.INIT_2E = INIT_2E;
defparam sb_ram8192x2r_inst.INIT_2F = INIT_2F;

defparam sb_ram8192x2r_inst.INIT_30 = INIT_30;
defparam sb_ram8192x2r_inst.INIT_31 = INIT_31;
defparam sb_ram8192x2r_inst.INIT_32 = INIT_32;
defparam sb_ram8192x2r_inst.INIT_33 = INIT_33;
defparam sb_ram8192x2r_inst.INIT_34 = INIT_34;
defparam sb_ram8192x2r_inst.INIT_35 = INIT_35;
defparam sb_ram8192x2r_inst.INIT_36 = INIT_36;
defparam sb_ram8192x2r_inst.INIT_37 = INIT_37;
defparam sb_ram8192x2r_inst.INIT_38 = INIT_38;
defparam sb_ram8192x2r_inst.INIT_39 = INIT_39;
defparam sb_ram8192x2r_inst.INIT_3A = INIT_3A;
defparam sb_ram8192x2r_inst.INIT_3B = INIT_3B;
defparam sb_ram8192x2r_inst.INIT_3C = INIT_3C;
defparam sb_ram8192x2r_inst.INIT_3D = INIT_3D;
defparam sb_ram8192x2r_inst.INIT_3E = INIT_3E;
defparam sb_ram8192x2r_inst.INIT_3F = INIT_3F;


`ifdef TIMINGCHECK
specify
   (RCLKN *> RDATA[0]) = (1.0, 1.0);
   (RCLKN *> RDATA[1]) = (1.0, 1.0);
   $setup(posedge WADDR[0], posedge WCLK, 1.0);
   $setup(negedge WADDR[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[0], 1.0);
   $hold(posedge WCLK, negedge WADDR[0], 1.0);
   $setup(posedge WADDR[1], posedge WCLK, 1.0);
   $setup(negedge WADDR[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[1], 1.0);
   $hold(posedge WCLK, negedge WADDR[1], 1.0);
   $setup(posedge WADDR[2], posedge WCLK, 1.0);
   $setup(negedge WADDR[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[2], 1.0);
   $hold(posedge WCLK, negedge WADDR[2], 1.0);
   $setup(posedge WADDR[3], posedge WCLK, 1.0);
   $setup(negedge WADDR[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[3], 1.0);
   $hold(posedge WCLK, negedge WADDR[3], 1.0);
   $setup(posedge WADDR[4], posedge WCLK, 1.0);
   $setup(negedge WADDR[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[4], 1.0);
   $hold(posedge WCLK, negedge WADDR[4], 1.0);
   $setup(posedge WADDR[5], posedge WCLK, 1.0);
   $setup(negedge WADDR[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[5], 1.0);
   $hold(posedge WCLK, negedge WADDR[5], 1.0);
   $setup(posedge WADDR[6], posedge WCLK, 1.0);
   $setup(negedge WADDR[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[6], 1.0);
   $hold(posedge WCLK, negedge WADDR[6], 1.0);
   $setup(posedge WADDR[7], posedge WCLK, 1.0);
   $setup(negedge WADDR[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[7], 1.0);
   $hold(posedge WCLK, negedge WADDR[7], 1.0);
   $setup(posedge WADDR[8], posedge WCLK, 1.0);
   $setup(negedge WADDR[8], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[8], 1.0);
   $hold(posedge WCLK, negedge WADDR[8], 1.0);
   $setup(posedge WADDR[9], posedge WCLK, 1.0);
   $setup(negedge WADDR[9], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[9], 1.0);
   $hold(posedge WCLK, negedge WADDR[9], 1.0);
   $setup(posedge WADDR[10], posedge WCLK, 1.0);
   $setup(negedge WADDR[10], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[10], 1.0);
   $hold(posedge WCLK, negedge WADDR[10], 1.0);
   $setup(posedge WADDR[11], posedge WCLK, 1.0);
   $setup(negedge WADDR[11], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[11], 1.0);
   $hold(posedge WCLK, negedge WADDR[11], 1.0);
   $setup(posedge WADDR[12], posedge WCLK, 1.0);
   $setup(negedge WADDR[12], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[12], 1.0);
   $hold(posedge WCLK, negedge WADDR[12], 1.0);
   $setup(posedge WDATA[0], posedge WCLK, 1.0);
   $setup(negedge WDATA[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[0], 1.0);
   $hold(posedge WCLK, negedge WDATA[0], 1.0);
   $setup(posedge WDATA[1], posedge WCLK, 1.0);
   $setup(negedge WDATA[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[1], 1.0);
   $hold(posedge WCLK, negedge WDATA[1], 1.0);
   $setup(posedge WCLKE, posedge WCLK, 1.0);
   $setup(negedge WCLKE, posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WCLKE, 1.0);
   $hold(posedge WCLK, negedge WCLKE, 1.0);
   $setup(posedge WE, posedge WCLK, 1.0);
   $setup(negedge WE, posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WE, 1.0);
   $hold(posedge WCLK, negedge WE, 1.0);
   $setup(posedge RADDR[0], posedge RCLKN, 1.0);
   $setup(negedge RADDR[0], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[0], 1.0);
   $hold(posedge RCLKN, negedge RADDR[0], 1.0);
   $setup(posedge RADDR[1], posedge RCLKN, 1.0);
   $setup(negedge RADDR[1], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[1], 1.0);
   $hold(posedge RCLKN, negedge RADDR[1], 1.0);
   $setup(posedge RADDR[2], posedge RCLKN, 1.0);
   $setup(negedge RADDR[2], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[2], 1.0);
   $hold(posedge RCLKN, negedge RADDR[2], 1.0);
   $setup(posedge RADDR[3], posedge RCLKN, 1.0);
   $setup(negedge RADDR[3], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[3], 1.0);
   $hold(posedge RCLKN, negedge RADDR[3], 1.0);
   $setup(posedge RADDR[4], posedge RCLKN, 1.0);
   $setup(negedge RADDR[4], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[4], 1.0);
   $hold(posedge RCLKN, negedge RADDR[4], 1.0);
   $setup(posedge RADDR[5], posedge RCLKN, 1.0);
   $setup(negedge RADDR[5], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[5], 1.0);
   $hold(posedge RCLKN, negedge RADDR[5], 1.0);
   $setup(posedge RADDR[6], posedge RCLKN, 1.0);
   $setup(negedge RADDR[6], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[6], 1.0);
   $hold(posedge RCLKN, negedge RADDR[6], 1.0);
   $setup(posedge RADDR[7], posedge RCLKN, 1.0);
   $setup(negedge RADDR[7], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[7], 1.0);
   $hold(posedge RCLKN, negedge RADDR[7], 1.0);
   $setup(posedge RADDR[8], posedge RCLKN, 1.0);
   $setup(negedge RADDR[8], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[8], 1.0);
   $hold(posedge RCLKN, negedge RADDR[8], 1.0);
   $setup(posedge RADDR[9], posedge RCLKN, 1.0);
   $setup(negedge RADDR[9], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[9], 1.0);
   $hold(posedge RCLKN, negedge RADDR[9], 1.0);
   $setup(posedge RADDR[10], posedge RCLKN, 1.0);
   $setup(negedge RADDR[10], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[10], 1.0);
   $hold(posedge RCLKN, negedge RADDR[10], 1.0);
   $setup(posedge RADDR[11], posedge RCLKN, 1.0);
   $setup(negedge RADDR[11], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[11], 1.0);
   $hold(posedge RCLKN, negedge RADDR[11], 1.0);
   $setup(posedge RADDR[12], posedge RCLKN, 1.0);
   $setup(negedge RADDR[12], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[12], 1.0);
   $hold(posedge RCLKN, negedge RADDR[12], 1.0);
   $setup(posedge RCLKE, posedge RCLKN, 1.0);
   $setup(negedge RCLKE, posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RCLKE, 1.0);
   $hold(posedge RCLKN, negedge RCLKE, 1.0);
   $setup(posedge RE, posedge RCLKN, 1.0);
   $setup(negedge RE, posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RE, 1.0);
   $hold(posedge RCLKN, negedge RE, 1.0);
endspecify
`endif

endmodule  // SB_RAM8192x2NR

//---------------------------------------
//	--- SB_RAM8192x2NW
//---------------------------------------
`timescale 1ps/1ps
module SB_RAM8192x2NW  ( RDATA, RCLK, RCLKE, RE, RADDR, WCLKN, WCLKE, WE, WADDR, WDATA ) ; 

output	[1:0]	RDATA;  
input         	RCLK;   
input           RCLKE; 
input           RE; 
input	[12:0]  RADDR; 
input           WCLKN; 
input           WCLKE; 
input           WE; 
input 	[12:0]  WADDR; 
input 	[1:0]	WDATA;  

parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;


wire WCLK;
assign (weak0, weak1) RCLKE =1'b1 ;
assign (weak0, weak1) RE =1'b0 ;
assign (weak0, weak1) WCLKE =1'b1 ;
assign (weak0, weak1) WE =1'b0 ;
assign WCLK = ~WCLKN;

SB_RAM8192x2 sb_ram8192x2w_inst (
	.RDATA(RDATA),
	.RCLK(RCLK),
	.RCLKE(RCLKE),
	.RE(RE),
	.RADDR(RADDR),
	.WCLK(WCLK),
	.WCLKE(WCLKE),
	.WE(WE),
	.WADDR(WADDR),
	.WDATA(WDATA));

defparam sb_ram8192x2w_inst.INIT_0 = INIT_0;
defparam sb_ram8192x2w_inst.INIT_1 = INIT_1;
defparam sb_ram8192x2w_inst.INIT_2 = INIT_2;
defparam sb_ram8192x2w_inst.INIT_3 = INIT_3;
defparam sb_ram8192x2w_inst.INIT_4 = INIT_4;
defparam sb_ram8192x2w_inst.INIT_5 = INIT_5;
defparam sb_ram8192x2w_inst.INIT_6 = INIT_6;
defparam sb_ram8192x2w_inst.INIT_7 = INIT_7;
defparam sb_ram8192x2w_inst.INIT_8 = INIT_8;
defparam sb_ram8192x2w_inst.INIT_9 = INIT_9;
defparam sb_ram8192x2w_inst.INIT_A = INIT_A;
defparam sb_ram8192x2w_inst.INIT_B = INIT_B;
defparam sb_ram8192x2w_inst.INIT_C = INIT_C;
defparam sb_ram8192x2w_inst.INIT_D = INIT_D;
defparam sb_ram8192x2w_inst.INIT_E = INIT_E;
defparam sb_ram8192x2w_inst.INIT_F = INIT_F;

defparam sb_ram8192x2w_inst.INIT_10 = INIT_10;
defparam sb_ram8192x2w_inst.INIT_11 = INIT_11;
defparam sb_ram8192x2w_inst.INIT_12 = INIT_12;
defparam sb_ram8192x2w_inst.INIT_13 = INIT_13;
defparam sb_ram8192x2w_inst.INIT_14 = INIT_14;
defparam sb_ram8192x2w_inst.INIT_15 = INIT_15;
defparam sb_ram8192x2w_inst.INIT_16 = INIT_16;
defparam sb_ram8192x2w_inst.INIT_17 = INIT_17;
defparam sb_ram8192x2w_inst.INIT_18 = INIT_18;
defparam sb_ram8192x2w_inst.INIT_19 = INIT_19;
defparam sb_ram8192x2w_inst.INIT_1A = INIT_1A;
defparam sb_ram8192x2w_inst.INIT_1B = INIT_1B;
defparam sb_ram8192x2w_inst.INIT_1C = INIT_1C;
defparam sb_ram8192x2w_inst.INIT_1D = INIT_1D;
defparam sb_ram8192x2w_inst.INIT_1E = INIT_1E;
defparam sb_ram8192x2w_inst.INIT_1F = INIT_1F;

defparam sb_ram8192x2w_inst.INIT_20 = INIT_20;
defparam sb_ram8192x2w_inst.INIT_21 = INIT_21;
defparam sb_ram8192x2w_inst.INIT_22 = INIT_22;
defparam sb_ram8192x2w_inst.INIT_23 = INIT_23;
defparam sb_ram8192x2w_inst.INIT_24 = INIT_24;
defparam sb_ram8192x2w_inst.INIT_25 = INIT_25;
defparam sb_ram8192x2w_inst.INIT_26 = INIT_26;
defparam sb_ram8192x2w_inst.INIT_27 = INIT_27;
defparam sb_ram8192x2w_inst.INIT_28 = INIT_28;
defparam sb_ram8192x2w_inst.INIT_29 = INIT_29;
defparam sb_ram8192x2w_inst.INIT_2A = INIT_2A;
defparam sb_ram8192x2w_inst.INIT_2B = INIT_2B;
defparam sb_ram8192x2w_inst.INIT_2C = INIT_2C;
defparam sb_ram8192x2w_inst.INIT_2D = INIT_2D;
defparam sb_ram8192x2w_inst.INIT_2E = INIT_2E;
defparam sb_ram8192x2w_inst.INIT_2F = INIT_2F;

defparam sb_ram8192x2w_inst.INIT_30 = INIT_30;
defparam sb_ram8192x2w_inst.INIT_31 = INIT_31;
defparam sb_ram8192x2w_inst.INIT_32 = INIT_32;
defparam sb_ram8192x2w_inst.INIT_33 = INIT_33;
defparam sb_ram8192x2w_inst.INIT_34 = INIT_34;
defparam sb_ram8192x2w_inst.INIT_35 = INIT_35;
defparam sb_ram8192x2w_inst.INIT_36 = INIT_36;
defparam sb_ram8192x2w_inst.INIT_37 = INIT_37;
defparam sb_ram8192x2w_inst.INIT_38 = INIT_38;
defparam sb_ram8192x2w_inst.INIT_39 = INIT_39;
defparam sb_ram8192x2w_inst.INIT_3A = INIT_3A;
defparam sb_ram8192x2w_inst.INIT_3B = INIT_3B;
defparam sb_ram8192x2w_inst.INIT_3C = INIT_3C;
defparam sb_ram8192x2w_inst.INIT_3D = INIT_3D;
defparam sb_ram8192x2w_inst.INIT_3E = INIT_3E;
defparam sb_ram8192x2w_inst.INIT_3F = INIT_3F;

`ifdef TIMINGCHECK
specify
   (RCLK *> RDATA[0]) = (1.0, 1.0);
   (RCLK *> RDATA[1]) = (1.0, 1.0);
   $setup(posedge WADDR[0], posedge WCLKN, 1.0);
   $setup(negedge WADDR[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[0], 1.0);
   $hold(posedge WCLKN, negedge WADDR[0], 1.0);
   $setup(posedge WADDR[1], posedge WCLKN, 1.0);
   $setup(negedge WADDR[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[1], 1.0);
   $hold(posedge WCLKN, negedge WADDR[1], 1.0);
   $setup(posedge WADDR[2], posedge WCLKN, 1.0);
   $setup(negedge WADDR[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[2], 1.0);
   $hold(posedge WCLKN, negedge WADDR[2], 1.0);
   $setup(posedge WADDR[3], posedge WCLKN, 1.0);
   $setup(negedge WADDR[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[3], 1.0);
   $hold(posedge WCLKN, negedge WADDR[3], 1.0);
   $setup(posedge WADDR[4], posedge WCLKN, 1.0);
   $setup(negedge WADDR[4], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[4], 1.0);
   $hold(posedge WCLKN, negedge WADDR[4], 1.0);
   $setup(posedge WADDR[5], posedge WCLKN, 1.0);
   $setup(negedge WADDR[5], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[5], 1.0);
   $hold(posedge WCLKN, negedge WADDR[5], 1.0);
   $setup(posedge WADDR[6], posedge WCLKN, 1.0);
   $setup(negedge WADDR[6], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[6], 1.0);
   $hold(posedge WCLKN, negedge WADDR[6], 1.0);
   $setup(posedge WADDR[7], posedge WCLKN, 1.0);
   $setup(negedge WADDR[7], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[7], 1.0);
   $hold(posedge WCLKN, negedge WADDR[7], 1.0);
   $setup(posedge WADDR[8], posedge WCLKN, 1.0);
   $setup(negedge WADDR[8], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[8], 1.0);
   $hold(posedge WCLKN, negedge WADDR[8], 1.0);
   $setup(posedge WADDR[9], posedge WCLKN, 1.0);
   $setup(negedge WADDR[9], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[9], 1.0);
   $hold(posedge WCLKN, negedge WADDR[9], 1.0);
   $setup(posedge WADDR[10], posedge WCLKN, 1.0);
   $setup(negedge WADDR[10], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[10], 1.0);
   $hold(posedge WCLKN, negedge WADDR[10], 1.0);
   $setup(posedge WADDR[11], posedge WCLKN, 1.0);
   $setup(negedge WADDR[11], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[11], 1.0);
   $hold(posedge WCLKN, negedge WADDR[11], 1.0);
   $setup(posedge WADDR[12], posedge WCLKN, 1.0);
   $setup(negedge WADDR[12], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[12], 1.0);
   $hold(posedge WCLKN, negedge WADDR[12], 1.0);
   $setup(posedge WDATA[0], posedge WCLKN, 1.0);
   $setup(negedge WDATA[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[0], 1.0);
   $hold(posedge WCLKN, negedge WDATA[0], 1.0);
   $setup(posedge WDATA[1], posedge WCLKN, 1.0);
   $setup(negedge WDATA[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[1], 1.0);
   $hold(posedge WCLKN, negedge WDATA[1], 1.0);
   $setup(posedge WCLKE, posedge WCLKN, 1.0);
   $setup(negedge WCLKE, posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WCLKE, 1.0);
   $hold(posedge WCLKN, negedge WCLKE, 1.0);
   $setup(posedge WE, posedge WCLKN, 1.0);
   $setup(negedge WE, posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WE, 1.0);
   $hold(posedge WCLKN, negedge WE, 1.0);
   $setup(posedge RADDR[0], posedge RCLK, 1.0);
   $setup(negedge RADDR[0], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[0], 1.0);
   $hold(posedge RCLK, negedge RADDR[0], 1.0);
   $setup(posedge RADDR[1], posedge RCLK, 1.0);
   $setup(negedge RADDR[1], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[1], 1.0);
   $hold(posedge RCLK, negedge RADDR[1], 1.0);
   $setup(posedge RADDR[2], posedge RCLK, 1.0);
   $setup(negedge RADDR[2], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[2], 1.0);
   $hold(posedge RCLK, negedge RADDR[2], 1.0);
   $setup(posedge RADDR[3], posedge RCLK, 1.0);
   $setup(negedge RADDR[3], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[3], 1.0);
   $hold(posedge RCLK, negedge RADDR[3], 1.0);
   $setup(posedge RADDR[4], posedge RCLK, 1.0);
   $setup(negedge RADDR[4], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[4], 1.0);
   $hold(posedge RCLK, negedge RADDR[4], 1.0);
   $setup(posedge RADDR[5], posedge RCLK, 1.0);
   $setup(negedge RADDR[5], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[5], 1.0);
   $hold(posedge RCLK, negedge RADDR[5], 1.0);
   $setup(posedge RADDR[6], posedge RCLK, 1.0);
   $setup(negedge RADDR[6], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[6], 1.0);
   $hold(posedge RCLK, negedge RADDR[6], 1.0);
   $setup(posedge RADDR[7], posedge RCLK, 1.0);
   $setup(negedge RADDR[7], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[7], 1.0);
   $hold(posedge RCLK, negedge RADDR[7], 1.0);
   $setup(posedge RADDR[8], posedge RCLK, 1.0);
   $setup(negedge RADDR[8], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[8], 1.0);
   $hold(posedge RCLK, negedge RADDR[8], 1.0);
   $setup(posedge RADDR[9], posedge RCLK, 1.0);
   $setup(negedge RADDR[9], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[9], 1.0);
   $hold(posedge RCLK, negedge RADDR[9], 1.0);
   $setup(posedge RADDR[10], posedge RCLK, 1.0);
   $setup(negedge RADDR[10], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[10], 1.0);
   $hold(posedge RCLK, negedge RADDR[10], 1.0);
   $setup(posedge RADDR[11], posedge RCLK, 1.0);
   $setup(negedge RADDR[11], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[11], 1.0);
   $hold(posedge RCLK, negedge RADDR[11], 1.0);
   $setup(posedge RADDR[12], posedge RCLK, 1.0);
   $setup(negedge RADDR[12], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[12], 1.0);
   $hold(posedge RCLK, negedge RADDR[12], 1.0);
   $setup(posedge RCLKE, posedge RCLK, 1.0);
   $setup(negedge RCLKE, posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RCLKE, 1.0);
   $hold(posedge RCLK, negedge RCLKE, 1.0);
   $setup(posedge RE, posedge RCLK, 1.0);
   $setup(negedge RE, posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RE, 1.0);
   $hold(posedge RCLK, negedge RE, 1.0);
endspecify
`endif

endmodule // SB_RAM8192x2NW 

//---------------------------------------
//	--- SB_RAM8192x2NRNW
//---------------------------------------
`timescale 1ps/1ps
module  SB_RAM8192x2NRNW  ( RDATA, RCLKN, RCLKE, RE, RADDR, WCLKN, WCLKE, WE, WADDR, WDATA ); 

output	[1:0]	RDATA;  
input         	RCLKN;   
input           RCLKE; 
input           RE; 
input	[12:0]  RADDR; 
input           WCLKN; 
input           WCLKE; 
input           WE; 
input 	[12:0]  WADDR; 
input 	[1:0]	WDATA; 

parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;


wire RCLK, WCLK;
assign (weak0, weak1) RCLKE =1'b1 ;
assign (weak0, weak1) RE =1'b0 ;
assign (weak0, weak1) WCLKE =1'b1 ;
assign (weak0, weak1) WE =1'b0 ;
assign RCLK = ~RCLKN;
assign WCLK = ~WCLKN;

SB_RAM8192x2 sb_ram8192x2rw_inst (
	.RDATA(RDATA),
	.RCLK(RCLK),
	.RCLKE(RCLKE),
	.RE(RE),
	.RADDR(RADDR),
	.WCLK(WCLK),
	.WCLKE(WCLKE),
	.WE(WE),
	.WADDR(WADDR),
	.WDATA(WDATA));

defparam sb_ram8192x2rw_inst.INIT_0 = INIT_0;
defparam sb_ram8192x2rw_inst.INIT_1 = INIT_1;
defparam sb_ram8192x2rw_inst.INIT_2 = INIT_2;
defparam sb_ram8192x2rw_inst.INIT_3 = INIT_3;
defparam sb_ram8192x2rw_inst.INIT_4 = INIT_4;
defparam sb_ram8192x2rw_inst.INIT_5 = INIT_5;
defparam sb_ram8192x2rw_inst.INIT_6 = INIT_6;
defparam sb_ram8192x2rw_inst.INIT_7 = INIT_7;
defparam sb_ram8192x2rw_inst.INIT_8 = INIT_8;
defparam sb_ram8192x2rw_inst.INIT_9 = INIT_9;
defparam sb_ram8192x2rw_inst.INIT_A = INIT_A;
defparam sb_ram8192x2rw_inst.INIT_B = INIT_B;
defparam sb_ram8192x2rw_inst.INIT_C = INIT_C;
defparam sb_ram8192x2rw_inst.INIT_D = INIT_D;
defparam sb_ram8192x2rw_inst.INIT_E = INIT_E;
defparam sb_ram8192x2rw_inst.INIT_F = INIT_F;

defparam sb_ram8192x2rw_inst.INIT_10 = INIT_10;
defparam sb_ram8192x2rw_inst.INIT_11 = INIT_11;
defparam sb_ram8192x2rw_inst.INIT_12 = INIT_12;
defparam sb_ram8192x2rw_inst.INIT_13 = INIT_13;
defparam sb_ram8192x2rw_inst.INIT_14 = INIT_14;
defparam sb_ram8192x2rw_inst.INIT_15 = INIT_15;
defparam sb_ram8192x2rw_inst.INIT_16 = INIT_16;
defparam sb_ram8192x2rw_inst.INIT_17 = INIT_17;
defparam sb_ram8192x2rw_inst.INIT_18 = INIT_18;
defparam sb_ram8192x2rw_inst.INIT_19 = INIT_19;
defparam sb_ram8192x2rw_inst.INIT_1A = INIT_1A;
defparam sb_ram8192x2rw_inst.INIT_1B = INIT_1B;
defparam sb_ram8192x2rw_inst.INIT_1C = INIT_1C;
defparam sb_ram8192x2rw_inst.INIT_1D = INIT_1D;
defparam sb_ram8192x2rw_inst.INIT_1E = INIT_1E;
defparam sb_ram8192x2rw_inst.INIT_1F = INIT_1F;

defparam sb_ram8192x2rw_inst.INIT_20 = INIT_20;
defparam sb_ram8192x2rw_inst.INIT_21 = INIT_21;
defparam sb_ram8192x2rw_inst.INIT_22 = INIT_22;
defparam sb_ram8192x2rw_inst.INIT_23 = INIT_23;
defparam sb_ram8192x2rw_inst.INIT_24 = INIT_24;
defparam sb_ram8192x2rw_inst.INIT_25 = INIT_25;
defparam sb_ram8192x2rw_inst.INIT_26 = INIT_26;
defparam sb_ram8192x2rw_inst.INIT_27 = INIT_27;
defparam sb_ram8192x2rw_inst.INIT_28 = INIT_28;
defparam sb_ram8192x2rw_inst.INIT_29 = INIT_29;
defparam sb_ram8192x2rw_inst.INIT_2A = INIT_2A;
defparam sb_ram8192x2rw_inst.INIT_2B = INIT_2B;
defparam sb_ram8192x2rw_inst.INIT_2C = INIT_2C;
defparam sb_ram8192x2rw_inst.INIT_2D = INIT_2D;
defparam sb_ram8192x2rw_inst.INIT_2E = INIT_2E;
defparam sb_ram8192x2rw_inst.INIT_2F = INIT_2F;

defparam sb_ram8192x2rw_inst.INIT_30 = INIT_30;
defparam sb_ram8192x2rw_inst.INIT_31 = INIT_31;
defparam sb_ram8192x2rw_inst.INIT_32 = INIT_32;
defparam sb_ram8192x2rw_inst.INIT_33 = INIT_33;
defparam sb_ram8192x2rw_inst.INIT_34 = INIT_34;
defparam sb_ram8192x2rw_inst.INIT_35 = INIT_35;
defparam sb_ram8192x2rw_inst.INIT_36 = INIT_36;
defparam sb_ram8192x2rw_inst.INIT_37 = INIT_37;
defparam sb_ram8192x2rw_inst.INIT_38 = INIT_38;
defparam sb_ram8192x2rw_inst.INIT_39 = INIT_39;
defparam sb_ram8192x2rw_inst.INIT_3A = INIT_3A;
defparam sb_ram8192x2rw_inst.INIT_3B = INIT_3B;
defparam sb_ram8192x2rw_inst.INIT_3C = INIT_3C;
defparam sb_ram8192x2rw_inst.INIT_3D = INIT_3D;
defparam sb_ram8192x2rw_inst.INIT_3E = INIT_3E;
defparam sb_ram8192x2rw_inst.INIT_3F = INIT_3F;


`ifdef TIMINGCHECK
specify
   (RCLKN *> RDATA[0]) = (1.0, 1.0);
   (RCLKN *> RDATA[1]) = (1.0, 1.0);
   $setup(posedge WADDR[0], posedge WCLKN, 1.0);
   $setup(negedge WADDR[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[0], 1.0);
   $hold(posedge WCLKN, negedge WADDR[0], 1.0);
   $setup(posedge WADDR[1], posedge WCLKN, 1.0);
   $setup(negedge WADDR[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[1], 1.0);
   $hold(posedge WCLKN, negedge WADDR[1], 1.0);
   $setup(posedge WADDR[2], posedge WCLKN, 1.0);
   $setup(negedge WADDR[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[2], 1.0);
   $hold(posedge WCLKN, negedge WADDR[2], 1.0);
   $setup(posedge WADDR[3], posedge WCLKN, 1.0);
   $setup(negedge WADDR[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[3], 1.0);
   $hold(posedge WCLKN, negedge WADDR[3], 1.0);
   $setup(posedge WADDR[4], posedge WCLKN, 1.0);
   $setup(negedge WADDR[4], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[4], 1.0);
   $hold(posedge WCLKN, negedge WADDR[4], 1.0);
   $setup(posedge WADDR[5], posedge WCLKN, 1.0);
   $setup(negedge WADDR[5], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[5], 1.0);
   $hold(posedge WCLKN, negedge WADDR[5], 1.0);
   $setup(posedge WADDR[6], posedge WCLKN, 1.0);
   $setup(negedge WADDR[6], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[6], 1.0);
   $hold(posedge WCLKN, negedge WADDR[6], 1.0);
   $setup(posedge WADDR[7], posedge WCLKN, 1.0);
   $setup(negedge WADDR[7], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[7], 1.0);
   $hold(posedge WCLKN, negedge WADDR[7], 1.0);
   $setup(posedge WADDR[8], posedge WCLKN, 1.0);
   $setup(negedge WADDR[8], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[8], 1.0);
   $hold(posedge WCLKN, negedge WADDR[8], 1.0);
   $setup(posedge WADDR[9], posedge WCLKN, 1.0);
   $setup(negedge WADDR[9], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[9], 1.0);
   $hold(posedge WCLKN, negedge WADDR[9], 1.0);
   $setup(posedge WADDR[10], posedge WCLKN, 1.0);
   $setup(negedge WADDR[10], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[10], 1.0);
   $hold(posedge WCLKN, negedge WADDR[10], 1.0);
   $setup(posedge WADDR[11], posedge WCLKN, 1.0);
   $setup(negedge WADDR[11], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[11], 1.0);
   $hold(posedge WCLKN, negedge WADDR[11], 1.0);
   $setup(posedge WADDR[12], posedge WCLKN, 1.0);
   $setup(negedge WADDR[12], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[12], 1.0);
   $hold(posedge WCLKN, negedge WADDR[12], 1.0);
   $setup(posedge WDATA[0], posedge WCLKN, 1.0);
   $setup(negedge WDATA[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[0], 1.0);
   $hold(posedge WCLKN, negedge WDATA[0], 1.0);
   $setup(posedge WDATA[1], posedge WCLKN, 1.0);
   $setup(negedge WDATA[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[1], 1.0);
   $hold(posedge WCLKN, negedge WDATA[1], 1.0);
   $setup(posedge WCLKE, posedge WCLKN, 1.0);
   $setup(negedge WCLKE, posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WCLKE, 1.0);
   $hold(posedge WCLKN, negedge WCLKE, 1.0);
   $setup(posedge WE, posedge WCLKN, 1.0);
   $setup(negedge WE, posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WE, 1.0);
   $hold(posedge WCLKN, negedge WE, 1.0);
   $setup(posedge RADDR[0], posedge RCLKN, 1.0);
   $setup(negedge RADDR[0], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[0], 1.0);
   $hold(posedge RCLKN, negedge RADDR[0], 1.0);
   $setup(posedge RADDR[1], posedge RCLKN, 1.0);
   $setup(negedge RADDR[1], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[1], 1.0);
   $hold(posedge RCLKN, negedge RADDR[1], 1.0);
   $setup(posedge RADDR[2], posedge RCLKN, 1.0);
   $setup(negedge RADDR[2], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[2], 1.0);
   $hold(posedge RCLKN, negedge RADDR[2], 1.0);
   $setup(posedge RADDR[3], posedge RCLKN, 1.0);
   $setup(negedge RADDR[3], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[3], 1.0);
   $hold(posedge RCLKN, negedge RADDR[3], 1.0);
   $setup(posedge RADDR[4], posedge RCLKN, 1.0);
   $setup(negedge RADDR[4], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[4], 1.0);
   $hold(posedge RCLKN, negedge RADDR[4], 1.0);
   $setup(posedge RADDR[5], posedge RCLKN, 1.0);
   $setup(negedge RADDR[5], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[5], 1.0);
   $hold(posedge RCLKN, negedge RADDR[5], 1.0);
   $setup(posedge RADDR[6], posedge RCLKN, 1.0);
   $setup(negedge RADDR[6], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[6], 1.0);
   $hold(posedge RCLKN, negedge RADDR[6], 1.0);
   $setup(posedge RADDR[7], posedge RCLKN, 1.0);
   $setup(negedge RADDR[7], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[7], 1.0);
   $hold(posedge RCLKN, negedge RADDR[7], 1.0);
   $setup(posedge RADDR[8], posedge RCLKN, 1.0);
   $setup(negedge RADDR[8], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[8], 1.0);
   $hold(posedge RCLKN, negedge RADDR[8], 1.0);
   $setup(posedge RADDR[9], posedge RCLKN, 1.0);
   $setup(negedge RADDR[9], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[9], 1.0);
   $hold(posedge RCLKN, negedge RADDR[9], 1.0);
   $setup(posedge RADDR[10], posedge RCLKN, 1.0);
   $setup(negedge RADDR[10], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[10], 1.0);
   $hold(posedge RCLKN, negedge RADDR[10], 1.0);
   $setup(posedge RADDR[11], posedge RCLKN, 1.0);
   $setup(negedge RADDR[11], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[11], 1.0);
   $hold(posedge RCLKN, negedge RADDR[11], 1.0);
   $setup(posedge RADDR[12], posedge RCLKN, 1.0);
   $setup(negedge RADDR[12], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[12], 1.0);
   $hold(posedge RCLKN, negedge RADDR[12], 1.0);
   $setup(posedge RCLKE, posedge RCLKN, 1.0);
   $setup(negedge RCLKE, posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RCLKE, 1.0);
   $hold(posedge RCLKN, negedge RCLKE, 1.0);
   $setup(posedge RE, posedge RCLKN, 1.0);
   $setup(negedge RE, posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RE, 1.0);
   $hold(posedge RCLKN, negedge RE, 1.0);
endspecify
`endif

endmodule // SB_RAM8192x2NRNW 

//---------------------------------------------------------------
//	 SB_RAM16K LeafLevel RamBlock for Physical Ram Wrappers      
//---------------------------------------------------------------
`timescale 1ps/1ps
module SB_RAM16K (RDATA, RCLK, RCLKE, RE, RADDR, WCLK, WCLKE, WE, WADDR, MASK, WDATA);
output [15:0] RDATA;
input RCLK;
input RCLKE;
input RE;
input [9:0] RADDR;
input WCLK;
input WCLKE;
input WE;
input [9:0] WADDR;
input [15:0] MASK;
input [15:0] WDATA;

parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

// local Parameters
localparam			CLOCK_PERIOD = 200;	//
localparam 			DELAY	= (CLOCK_PERIOD/10);		// Clock-to-output delay. Zero
							// time delays can be confusing
							// and sometimes cause problems.
localparam 			BUS_WIDTH = 16;		// Width of RAM (number of bits)

localparam 			ADDRESS_BUS_SIZE = 10;	// Number of bits required to
							// represent the RAM address

localparam   ADDRESSABLE_SPACE  = 2**ADDRESS_BUS_SIZE;	// Decimal address range [2^Size:0]


// SIGNAL DECLARATIONS
wire			   	WCLK_g, RCLK_g;
reg 				WCLKE_sync, RCLKE_sync; 
assign (weak0, weak1) RCLKE =1'b1 ;
assign (weak0, weak1) RE =1'b0 ;
assign (weak0, weak1) WCLKE =1'b1 ;
assign (weak0, weak1) WE =1'b0 ;

assign (weak0, weak1) MASK = 16'b0;

//reg  [BUS_WIDTH-1:0] Memory [ADDRESSABLE_SPACE-1:0];	// The RAM
reg	Memory	[BUS_WIDTH*ADDRESSABLE_SPACE-1:0];
// 
event Read_e, Write_e;

//////////////////// Collision detect begins here ///////////////////////////////
localparam 	TRUE = 1'b1;
localparam	FALSE = 1'b0;
reg 		Time_Collision_Detected = 1'b0;
wire		Address_Collision_Detected;

event Collision_e;

time COLLISION_TIME_WINDOW = (CLOCK_PERIOD/8); // This is an arbitray value, but is better than using an absolute 
						    // value, because the actual time window depends on the actual silicon 
						    // implementation. Thus the test is indicative of an Error and not
						    // guaranteed to be an error. Even so this is usefull.
time time_WCLK_RCLK, time_WCLK, time_RCLK;


//function reg Check_Timed_Window_Violation;
function	Check_Timed_Window_Violation;	//	by Jeffrey
input T1, T2, Minimum_Time_Window;
time T1, T2;
time Minimum_Time_Window;
time Difference;	
	begin
		Difference = (T1 - T2);
		if (Difference < 0) Difference = -Difference;
		Check_Timed_Window_Violation = (Difference < Minimum_Time_Window);
	end
endfunction


initial begin
       time_WCLK = CLOCK_PERIOD;	// Arbitrary initialisation value, ensure no window collison error on first clock edge.
       time_RCLK = (CLOCK_PERIOD*8);	// Arbitrary initialisation difference value, ensure no collision error on first clock edge.					
end

integer	i,j;

genvar k;
wire [9:0] RADDR_g;
wire [9:0] WADDR_g;
wire [15:0] WDATA_g;
for (k = 0; k < 10; k = k + 1) begin
	assign RADDR_g[k] = (RADDR[k] === 1'bz)? 1'b0 : RADDR[k];
	assign WADDR_g[k] = (WADDR[k] === 1'bz)? 1'b0 : WADDR[k];
	assign WDATA_g[k] = (WDATA[k] === 1'bz)? 1'b0 : WDATA[k];
	assign WDATA_g[k+6] = (WDATA[k+6] === 1'bz)? 1'b0 : WDATA[k+6];
end

initial	//	initialize ram16k by init parameters, section by section
begin
	for	(i=0; i<=256/BUS_WIDTH -1; i=i+1)
	begin
		for	(j=0; j<=BUS_WIDTH-1; j=j+1)
		begin 

			Memory[BUS_WIDTH*i+j]		=	INIT_0[BUS_WIDTH*i+j];
			Memory[256*1+BUS_WIDTH*i+j]	=	INIT_1[BUS_WIDTH*i+j];
			Memory[256*2+BUS_WIDTH*i+j]	=	INIT_2[BUS_WIDTH*i+j];
			Memory[256*3+BUS_WIDTH*i+j]	=	INIT_3[BUS_WIDTH*i+j];
			Memory[256*4+BUS_WIDTH*i+j]	=	INIT_4[BUS_WIDTH*i+j];
			Memory[256*5+BUS_WIDTH*i+j]	=	INIT_5[BUS_WIDTH*i+j];
			Memory[256*6+BUS_WIDTH*i+j]	=	INIT_6[BUS_WIDTH*i+j];
			Memory[256*7+BUS_WIDTH*i+j]	=	INIT_7[BUS_WIDTH*i+j];
			Memory[256*8+BUS_WIDTH*i+j]	=	INIT_8[BUS_WIDTH*i+j];
			Memory[256*9+BUS_WIDTH*i+j]	=	INIT_9[BUS_WIDTH*i+j];
			Memory[256*10+BUS_WIDTH*i+j]	=	INIT_A[BUS_WIDTH*i+j];
			Memory[256*11+BUS_WIDTH*i+j]	=	INIT_B[BUS_WIDTH*i+j];
			Memory[256*12+BUS_WIDTH*i+j]	=	INIT_C[BUS_WIDTH*i+j];
			Memory[256*13+BUS_WIDTH*i+j]	=	INIT_D[BUS_WIDTH*i+j];
			Memory[256*14+BUS_WIDTH*i+j]	=	INIT_E[BUS_WIDTH*i+j];
			Memory[256*15+BUS_WIDTH*i+j]	=	INIT_F[BUS_WIDTH*i+j];

			Memory[256*16+BUS_WIDTH*i+j]	=	INIT_10[BUS_WIDTH*i+j];
			Memory[256*17+BUS_WIDTH*i+j]	=	INIT_11[BUS_WIDTH*i+j];
			Memory[256*18+BUS_WIDTH*i+j]	=	INIT_12[BUS_WIDTH*i+j];
			Memory[256*19+BUS_WIDTH*i+j]	=	INIT_13[BUS_WIDTH*i+j];
			Memory[256*20+BUS_WIDTH*i+j]	=	INIT_14[BUS_WIDTH*i+j];
			Memory[256*21+BUS_WIDTH*i+j]	=	INIT_15[BUS_WIDTH*i+j];
			Memory[256*22+BUS_WIDTH*i+j]	=	INIT_16[BUS_WIDTH*i+j];
			Memory[256*23+BUS_WIDTH*i+j]	=	INIT_17[BUS_WIDTH*i+j];
			Memory[256*24+BUS_WIDTH*i+j]	=	INIT_18[BUS_WIDTH*i+j];
			Memory[256*25+BUS_WIDTH*i+j]	=	INIT_19[BUS_WIDTH*i+j];
			Memory[256*26+BUS_WIDTH*i+j]	=	INIT_1A[BUS_WIDTH*i+j];
			Memory[256*27+BUS_WIDTH*i+j]	=	INIT_1B[BUS_WIDTH*i+j];
			Memory[256*28+BUS_WIDTH*i+j]	=	INIT_1C[BUS_WIDTH*i+j];
			Memory[256*29+BUS_WIDTH*i+j]	=	INIT_1D[BUS_WIDTH*i+j];
			Memory[256*30+BUS_WIDTH*i+j]	=	INIT_1E[BUS_WIDTH*i+j];
			Memory[256*31+BUS_WIDTH*i+j]	=	INIT_1F[BUS_WIDTH*i+j];

			Memory[256*32+BUS_WIDTH*i+j]	=	INIT_20[BUS_WIDTH*i+j];
			Memory[256*33+BUS_WIDTH*i+j]	=	INIT_21[BUS_WIDTH*i+j];
			Memory[256*34+BUS_WIDTH*i+j]	=	INIT_22[BUS_WIDTH*i+j];
			Memory[256*35+BUS_WIDTH*i+j]	=	INIT_23[BUS_WIDTH*i+j];
			Memory[256*36+BUS_WIDTH*i+j]	=	INIT_24[BUS_WIDTH*i+j];
			Memory[256*37+BUS_WIDTH*i+j]	=	INIT_25[BUS_WIDTH*i+j];
			Memory[256*38+BUS_WIDTH*i+j]	=	INIT_26[BUS_WIDTH*i+j];
			Memory[256*39+BUS_WIDTH*i+j]	=	INIT_27[BUS_WIDTH*i+j];
			Memory[256*40+BUS_WIDTH*i+j]	=	INIT_28[BUS_WIDTH*i+j];
			Memory[256*41+BUS_WIDTH*i+j]	=	INIT_29[BUS_WIDTH*i+j];
			Memory[256*42+BUS_WIDTH*i+j]	=	INIT_2A[BUS_WIDTH*i+j];
			Memory[256*43+BUS_WIDTH*i+j]	=	INIT_2B[BUS_WIDTH*i+j];
			Memory[256*44+BUS_WIDTH*i+j]	=	INIT_2C[BUS_WIDTH*i+j];
			Memory[256*45+BUS_WIDTH*i+j]	=	INIT_2D[BUS_WIDTH*i+j];
			Memory[256*46+BUS_WIDTH*i+j]	=	INIT_2E[BUS_WIDTH*i+j];
			Memory[256*47+BUS_WIDTH*i+j]	=	INIT_2F[BUS_WIDTH*i+j];

			Memory[256*48+BUS_WIDTH*i+j]	=	INIT_30[BUS_WIDTH*i+j];
			Memory[256*49+BUS_WIDTH*i+j]	=	INIT_31[BUS_WIDTH*i+j];
			Memory[256*50+BUS_WIDTH*i+j]	=	INIT_32[BUS_WIDTH*i+j];
			Memory[256*51+BUS_WIDTH*i+j]	=	INIT_33[BUS_WIDTH*i+j];
			Memory[256*52+BUS_WIDTH*i+j]	=	INIT_34[BUS_WIDTH*i+j];
			Memory[256*53+BUS_WIDTH*i+j]	=	INIT_35[BUS_WIDTH*i+j];
			Memory[256*54+BUS_WIDTH*i+j]	=	INIT_36[BUS_WIDTH*i+j];
			Memory[256*55+BUS_WIDTH*i+j]	=	INIT_37[BUS_WIDTH*i+j];
			Memory[256*56+BUS_WIDTH*i+j]	=	INIT_38[BUS_WIDTH*i+j];
			Memory[256*57+BUS_WIDTH*i+j]	=	INIT_39[BUS_WIDTH*i+j];
			Memory[256*58+BUS_WIDTH*i+j]	=	INIT_3A[BUS_WIDTH*i+j];
			Memory[256*59+BUS_WIDTH*i+j]	=	INIT_3B[BUS_WIDTH*i+j];
			Memory[256*60+BUS_WIDTH*i+j]	=	INIT_3C[BUS_WIDTH*i+j];
			Memory[256*61+BUS_WIDTH*i+j]	=	INIT_3D[BUS_WIDTH*i+j];
			Memory[256*62+BUS_WIDTH*i+j]	=	INIT_3E[BUS_WIDTH*i+j];
			Memory[256*63+BUS_WIDTH*i+j]	=	INIT_3F[BUS_WIDTH*i+j];
		end 
	end
end

assign Address_Collision_Detected = ((RE & WE & WCLKE & RCLKE)&(WADDR == RADDR)); 

always @(WCLK or WCLKE) 
begin 
	if(~WCLK)
	WCLKE_sync = WCLKE;   	
end 

always @(RCLK or RCLKE) 
begin 
	if (~RCLK)
	RCLKE_sync = RCLKE; 	
end 

assign WCLK_g = WCLK & WCLKE_sync;
assign RCLK_g = RCLK & RCLKE_sync;

always @(posedge WCLK_g) begin
	time_WCLK = $time;
end

always @(posedge RCLK_g) begin
    	time_RCLK = $time;
end
integer	SB_RAM16K_RDATA_log_file;									//.....................
initial	SB_RAM16K_RDATA_log_file=("SB_RAM16K_RDATA_log_file.txt");	//.....................
always @(posedge WCLK_g) begin

	Time_Collision_Detected = Check_Timed_Window_Violation(time_WCLK,time_RCLK,COLLISION_TIME_WINDOW);
        if (Time_Collision_Detected & Address_Collision_Detected)begin
        	$display("Warning: Write-Read collision detected, Data read value is XXXX\n");
 		$display("WCLK Time: %.3f   RCLK Time:%.3f  ",time_WCLK, time_RCLK,"WADDR: %d   RADDR:%d\n",WADDR, RADDR); 
 		$fdisplay(SB_RAM16K_RDATA_log_file,"Warning: Write-Read collision detected, Data read value is XXXX\n");
		$fdisplay(SB_RAM16K_RDATA_log_file,"WCLK Time: %.3f   RCLK Time:%.3f  ",time_WCLK, time_RCLK, "WADDR: %d   RADDR:%d\n",WADDR, RADDR); 	
 		-> Collision_e;
	end
end

//	code modify for universal verilog compiler

always @ (posedge WCLK_g)
begin
	if	(WE)
	begin
		-> Write_e;
		for	(i=0;i<=BUS_WIDTH-1; i=i+1)
		begin
			if	(MASK[i] !=1)
				Memory[WADDR_g*BUS_WIDTH+i]	<=	WDATA_g[i];
			else
				Memory[WADDR_g*BUS_WIDTH+i]	<=	Memory[WADDR_g*BUS_WIDTH+i];
		end
	end
end

reg	[BUS_WIDTH-1:0]	RDATA = 0;

// Look at the rising edge of the clock

always @ (posedge RCLK_g)
begin
	if	(RE)
	begin
		-> Read_e;
		if	(Time_Collision_Detected & Address_Collision_Detected) 
			RDATA <= {BUS_WIDTH{1'hX}};
		else
			for	(i=0;i<=BUS_WIDTH-1;i=i+1)
				RDATA[i]	<= Memory[RADDR_g*BUS_WIDTH+i];
	end
end

`ifdef TIMINGCHECK
specify
   (RCLK *> RDATA[0]) = (1.0, 1.0);
   (RCLK *> RDATA[1]) = (1.0, 1.0);
   (RCLK *> RDATA[2]) = (1.0, 1.0);
   (RCLK *> RDATA[3]) = (1.0, 1.0);
   (RCLK *> RDATA[4]) = (1.0, 1.0);
   (RCLK *> RDATA[5]) = (1.0, 1.0);
   (RCLK *> RDATA[6]) = (1.0, 1.0);
   (RCLK *> RDATA[7]) = (1.0, 1.0);
   (RCLK *> RDATA[8]) = (1.0, 1.0);
   (RCLK *> RDATA[9]) = (1.0, 1.0);
   (RCLK *> RDATA[10]) = (1.0, 1.0);
   (RCLK *> RDATA[11]) = (1.0, 1.0);
   (RCLK *> RDATA[12]) = (1.0, 1.0);
   (RCLK *> RDATA[13]) = (1.0, 1.0);
   (RCLK *> RDATA[14]) = (1.0, 1.0);
   (RCLK *> RDATA[15]) = (1.0, 1.0);
   $setup(posedge MASK[0], posedge WCLK, 1.0);
   $setup(negedge MASK[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[0], 1.0);
   $hold(posedge WCLK, negedge MASK[0], 1.0);
   $setup(posedge MASK[1], posedge WCLK, 1.0);
   $setup(negedge MASK[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[1], 1.0);
   $hold(posedge WCLK, negedge MASK[1], 1.0);
   $setup(posedge MASK[2], posedge WCLK, 1.0);
   $setup(negedge MASK[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[2], 1.0);
   $hold(posedge WCLK, negedge MASK[2], 1.0);
   $setup(posedge MASK[3], posedge WCLK, 1.0);
   $setup(negedge MASK[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[3], 1.0);
   $hold(posedge WCLK, negedge MASK[3], 1.0);
   $setup(posedge MASK[4], posedge WCLK, 1.0);
   $setup(negedge MASK[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[4], 1.0);
   $hold(posedge WCLK, negedge MASK[4], 1.0);
   $setup(posedge MASK[5], posedge WCLK, 1.0);
   $setup(negedge MASK[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[5], 1.0);
   $hold(posedge WCLK, negedge MASK[5], 1.0);
   $setup(posedge MASK[6], posedge WCLK, 1.0);
   $setup(negedge MASK[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[6], 1.0);
   $hold(posedge WCLK, negedge MASK[6], 1.0);
   $setup(posedge MASK[7], posedge WCLK, 1.0);
   $setup(negedge MASK[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[7], 1.0);
   $hold(posedge WCLK, negedge MASK[7], 1.0);
   $setup(posedge MASK[8], posedge WCLK, 1.0);
   $setup(negedge MASK[8], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[8], 1.0);
   $hold(posedge WCLK, negedge MASK[8], 1.0);
   $setup(posedge MASK[9], posedge WCLK, 1.0);
   $setup(negedge MASK[9], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[9], 1.0);
   $hold(posedge WCLK, negedge MASK[9], 1.0);
   $setup(posedge MASK[10], posedge WCLK, 1.0);
   $setup(negedge MASK[10], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[10], 1.0);
   $hold(posedge WCLK, negedge MASK[10], 1.0);
   $setup(posedge MASK[11], posedge WCLK, 1.0);
   $setup(negedge MASK[11], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[11], 1.0);
   $hold(posedge WCLK, negedge MASK[11], 1.0);
   $setup(posedge MASK[12], posedge WCLK, 1.0);
   $setup(negedge MASK[12], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[12], 1.0);
   $hold(posedge WCLK, negedge MASK[12], 1.0);
   $setup(posedge MASK[13], posedge WCLK, 1.0);
   $setup(negedge MASK[13], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[13], 1.0);
   $hold(posedge WCLK, negedge MASK[13], 1.0);
   $setup(posedge MASK[14], posedge WCLK, 1.0);
   $setup(negedge MASK[14], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[14], 1.0);
   $hold(posedge WCLK, negedge MASK[14], 1.0);
   $setup(posedge MASK[15], posedge WCLK, 1.0);
   $setup(negedge MASK[15], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[15], 1.0);
   $hold(posedge WCLK, negedge MASK[15], 1.0);
   $setup(posedge WADDR[0], posedge WCLK, 1.0);
   $setup(negedge WADDR[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[0], 1.0);
   $hold(posedge WCLK, negedge WADDR[0], 1.0);
   $setup(posedge WADDR[1], posedge WCLK, 1.0);
   $setup(negedge WADDR[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[1], 1.0);
   $hold(posedge WCLK, negedge WADDR[1], 1.0);
   $setup(posedge WADDR[2], posedge WCLK, 1.0);
   $setup(negedge WADDR[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[2], 1.0);
   $hold(posedge WCLK, negedge WADDR[2], 1.0);
   $setup(posedge WADDR[3], posedge WCLK, 1.0);
   $setup(negedge WADDR[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[3], 1.0);
   $hold(posedge WCLK, negedge WADDR[3], 1.0);
   $setup(posedge WADDR[4], posedge WCLK, 1.0);
   $setup(negedge WADDR[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[4], 1.0);
   $hold(posedge WCLK, negedge WADDR[4], 1.0);
   $setup(posedge WADDR[5], posedge WCLK, 1.0);
   $setup(negedge WADDR[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[5], 1.0);
   $hold(posedge WCLK, negedge WADDR[5], 1.0);
   $setup(posedge WADDR[6], posedge WCLK, 1.0);
   $setup(negedge WADDR[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[6], 1.0);
   $hold(posedge WCLK, negedge WADDR[6], 1.0);
   $setup(posedge WADDR[7], posedge WCLK, 1.0);
   $setup(negedge WADDR[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[7], 1.0);
   $hold(posedge WCLK, negedge WADDR[7], 1.0);
   $setup(posedge WADDR[8], posedge WCLK, 1.0);
   $setup(negedge WADDR[8], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[8], 1.0);
   $hold(posedge WCLK, negedge WADDR[8], 1.0);
   $setup(posedge WADDR[9], posedge WCLK, 1.0);
   $setup(negedge WADDR[9], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[9], 1.0);
   $hold(posedge WCLK, negedge WADDR[9], 1.0);
   $setup(posedge WDATA[0], posedge WCLK, 1.0);
   $setup(negedge WDATA[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[0], 1.0);
   $hold(posedge WCLK, negedge WDATA[0], 1.0);
   $setup(posedge WDATA[1], posedge WCLK, 1.0);
   $setup(negedge WDATA[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[1], 1.0);
   $hold(posedge WCLK, negedge WDATA[1], 1.0);
   $setup(posedge WDATA[2], posedge WCLK, 1.0);
   $setup(negedge WDATA[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[2], 1.0);
   $hold(posedge WCLK, negedge WDATA[2], 1.0);
   $setup(posedge WDATA[3], posedge WCLK, 1.0);
   $setup(negedge WDATA[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[3], 1.0);
   $hold(posedge WCLK, negedge WDATA[3], 1.0);
   $setup(posedge WDATA[4], posedge WCLK, 1.0);
   $setup(negedge WDATA[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[4], 1.0);
   $hold(posedge WCLK, negedge WDATA[4], 1.0);
   $setup(posedge WDATA[5], posedge WCLK, 1.0);
   $setup(negedge WDATA[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[5], 1.0);
   $hold(posedge WCLK, negedge WDATA[5], 1.0);
   $setup(posedge WDATA[6], posedge WCLK, 1.0);
   $setup(negedge WDATA[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[6], 1.0);
   $hold(posedge WCLK, negedge WDATA[6], 1.0);
   $setup(posedge WDATA[7], posedge WCLK, 1.0);
   $setup(negedge WDATA[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[7], 1.0);
   $hold(posedge WCLK, negedge WDATA[7], 1.0);
   $setup(posedge WDATA[8], posedge WCLK, 1.0);
   $setup(negedge WDATA[8], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[8], 1.0);
   $hold(posedge WCLK, negedge WDATA[8], 1.0);
   $setup(posedge WDATA[9], posedge WCLK, 1.0);
   $setup(negedge WDATA[9], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[9], 1.0);
   $hold(posedge WCLK, negedge WDATA[9], 1.0);
   $setup(posedge WDATA[10], posedge WCLK, 1.0);
   $setup(negedge WDATA[10], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[10], 1.0);
   $hold(posedge WCLK, negedge WDATA[10], 1.0);
   $setup(posedge WDATA[11], posedge WCLK, 1.0);
   $setup(negedge WDATA[11], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[11], 1.0);
   $hold(posedge WCLK, negedge WDATA[11], 1.0);
   $setup(posedge WDATA[12], posedge WCLK, 1.0);
   $setup(negedge WDATA[12], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[12], 1.0);
   $hold(posedge WCLK, negedge WDATA[12], 1.0);
   $setup(posedge WDATA[13], posedge WCLK, 1.0);
   $setup(negedge WDATA[13], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[13], 1.0);
   $hold(posedge WCLK, negedge WDATA[13], 1.0);
   $setup(posedge WDATA[14], posedge WCLK, 1.0);
   $setup(negedge WDATA[14], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[14], 1.0);
   $hold(posedge WCLK, negedge WDATA[14], 1.0);
   $setup(posedge WDATA[15], posedge WCLK, 1.0);
   $setup(negedge WDATA[15], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[15], 1.0);
   $hold(posedge WCLK, negedge WDATA[15], 1.0);
   $setup(posedge WCLKE, posedge WCLK, 1.0);
   $setup(negedge WCLKE, posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WCLKE, 1.0);
   $hold(posedge WCLK, negedge WCLKE, 1.0);
   $setup(posedge WE, posedge WCLK, 1.0);
   $setup(negedge WE, posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WE, 1.0);
   $hold(posedge WCLK, negedge WE, 1.0);
   $setup(posedge RADDR[0], posedge RCLK, 1.0);
   $setup(negedge RADDR[0], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[0], 1.0);
   $hold(posedge RCLK, negedge RADDR[0], 1.0);
   $setup(posedge RADDR[1], posedge RCLK, 1.0);
   $setup(negedge RADDR[1], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[1], 1.0);
   $hold(posedge RCLK, negedge RADDR[1], 1.0);
   $setup(posedge RADDR[2], posedge RCLK, 1.0);
   $setup(negedge RADDR[2], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[2], 1.0);
   $hold(posedge RCLK, negedge RADDR[2], 1.0);
   $setup(posedge RADDR[3], posedge RCLK, 1.0);
   $setup(negedge RADDR[3], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[3], 1.0);
   $hold(posedge RCLK, negedge RADDR[3], 1.0);
   $setup(posedge RADDR[4], posedge RCLK, 1.0);
   $setup(negedge RADDR[4], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[4], 1.0);
   $hold(posedge RCLK, negedge RADDR[4], 1.0);
   $setup(posedge RADDR[5], posedge RCLK, 1.0);
   $setup(negedge RADDR[5], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[5], 1.0);
   $hold(posedge RCLK, negedge RADDR[5], 1.0);
   $setup(posedge RADDR[6], posedge RCLK, 1.0);
   $setup(negedge RADDR[6], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[6], 1.0);
   $hold(posedge RCLK, negedge RADDR[6], 1.0);
   $setup(posedge RADDR[7], posedge RCLK, 1.0);
   $setup(negedge RADDR[7], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[7], 1.0);
   $hold(posedge RCLK, negedge RADDR[7], 1.0);
   $setup(posedge RADDR[8], posedge RCLK, 1.0);
   $setup(negedge RADDR[8], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[8], 1.0);
   $hold(posedge RCLK, negedge RADDR[8], 1.0);
   $setup(posedge RADDR[9], posedge RCLK, 1.0);
   $setup(negedge RADDR[9], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[9], 1.0);
   $hold(posedge RCLK, negedge RADDR[9], 1.0);
   $setup(posedge RCLKE, posedge RCLK, 1.0);
   $setup(negedge RCLKE, posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RCLKE, 1.0);
   $hold(posedge RCLK, negedge RCLKE, 1.0);
   $setup(posedge RE, posedge RCLK, 1.0);
   $setup(negedge RE, posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RE, 1.0);
   $hold(posedge RCLK, negedge RE, 1.0);
endspecify
`endif

endmodule	 //	SB_RAM16K

//-------------------------------------------
//   --SB_RAM40_16K 
//------------------------------------------- 

`timescale 1ps/1ps
module SB_RAM40_16K ( RDATA, RCLK, RCLKE, RE, RADDR, WCLK, WCLKE, WE, WADDR, MASK, WDATA ); 

output	[15:0]	RDATA;  
input         	RCLK;   
input           RCLKE; 
input           RE; 
input	[12:0]  RADDR; 
input           WCLK; 
input           WCLKE; 
input           WE; 
input 	[12:0]  WADDR; 
input 	[15:0]  MASK; 
input 	[15:0]	WDATA; 


parameter WRITE_MODE = 0;    // Configure Write Port as 1024x16 (0)/ 20148x8 (1)/ 4096x4 (2)/ 8192x2 (3)     
parameter READ_MODE  = 0;    // Configure Read  Port as 1024x16 (0)/ 20148x8 (1)/ 4096x4 (2)/ 8192x2 (3)

parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;  
 

assign (weak0, weak1) MASK = 16'b0;

wire [15:0] RD;
wire [15:0] WD;
wire [15:0] MASK_RAM;

reg [12:10] RADDR_reg;
always @(posedge RCLK) begin
	RADDR_reg[12:10] <= RADDR[12:10];
end

read_data_decoder read_decoder_inst (
	.di(RD),
	.ai(RADDR_reg[12:10]),
	.do(RDATA)
);
defparam read_decoder_inst.READ_MODE = READ_MODE;

write_data_decoder write_decoder_inst (
	.di(WDATA),
	.do(WD)
);
defparam write_decoder_inst.WRITE_MODE = WRITE_MODE;

mask_decoder mask_decoder_inst(
	.mi(MASK),
	.ai(WADDR[12:10]),
	.mo(MASK_RAM)
);
defparam mask_decoder_inst.WRITE_MODE = WRITE_MODE;

SB_RAM16K ram_inst (
	.RDATA(RD),
	.RCLK(RCLK),
	.RCLKE(RCLKE),
	.RE(RE),
	.RADDR(RADDR[9:0]),
	.WCLK(WCLK),
	.WCLKE(WCLKE),
	.WE(WE),
	.WADDR(WADDR[9:0]),
	.MASK(MASK_RAM),
	.WDATA(WD));

defparam ram_inst.INIT_0 = INIT_0;
defparam ram_inst.INIT_1 = INIT_1;
defparam ram_inst.INIT_2 = INIT_2;
defparam ram_inst.INIT_3 = INIT_3;
defparam ram_inst.INIT_4 = INIT_4;
defparam ram_inst.INIT_5 = INIT_5;
defparam ram_inst.INIT_6 = INIT_6;
defparam ram_inst.INIT_7 = INIT_7;
defparam ram_inst.INIT_8 = INIT_8;
defparam ram_inst.INIT_9 = INIT_9;
defparam ram_inst.INIT_A = INIT_A;
defparam ram_inst.INIT_B = INIT_B;
defparam ram_inst.INIT_C = INIT_C;
defparam ram_inst.INIT_D = INIT_D;
defparam ram_inst.INIT_E = INIT_E;
defparam ram_inst.INIT_F = INIT_F;

defparam ram_inst.INIT_10 = INIT_10;
defparam ram_inst.INIT_11 = INIT_11;
defparam ram_inst.INIT_12 = INIT_12;
defparam ram_inst.INIT_13 = INIT_13;
defparam ram_inst.INIT_14 = INIT_14;
defparam ram_inst.INIT_15 = INIT_15;
defparam ram_inst.INIT_16 = INIT_16;
defparam ram_inst.INIT_17 = INIT_17;
defparam ram_inst.INIT_18 = INIT_18;
defparam ram_inst.INIT_19 = INIT_19;
defparam ram_inst.INIT_1A = INIT_1A;
defparam ram_inst.INIT_1B = INIT_1B;
defparam ram_inst.INIT_1C = INIT_1C;
defparam ram_inst.INIT_1D = INIT_1D;
defparam ram_inst.INIT_1E = INIT_1E;
defparam ram_inst.INIT_1F = INIT_1F;

defparam ram_inst.INIT_20 = INIT_20;
defparam ram_inst.INIT_21 = INIT_21;
defparam ram_inst.INIT_22 = INIT_22;
defparam ram_inst.INIT_23 = INIT_23;
defparam ram_inst.INIT_24 = INIT_24;
defparam ram_inst.INIT_25 = INIT_25;
defparam ram_inst.INIT_26 = INIT_26;
defparam ram_inst.INIT_27 = INIT_27;
defparam ram_inst.INIT_28 = INIT_28;
defparam ram_inst.INIT_29 = INIT_29;
defparam ram_inst.INIT_2A = INIT_2A;
defparam ram_inst.INIT_2B = INIT_2B;
defparam ram_inst.INIT_2C = INIT_2C;
defparam ram_inst.INIT_2D = INIT_2D;
defparam ram_inst.INIT_2E = INIT_2E;
defparam ram_inst.INIT_2F = INIT_2F;

defparam ram_inst.INIT_30 = INIT_30;
defparam ram_inst.INIT_31 = INIT_31;
defparam ram_inst.INIT_32 = INIT_32;
defparam ram_inst.INIT_33 = INIT_33;
defparam ram_inst.INIT_34 = INIT_34;
defparam ram_inst.INIT_35 = INIT_35;
defparam ram_inst.INIT_36 = INIT_36;
defparam ram_inst.INIT_37 = INIT_37;
defparam ram_inst.INIT_38 = INIT_38;
defparam ram_inst.INIT_39 = INIT_39;
defparam ram_inst.INIT_3A = INIT_3A;
defparam ram_inst.INIT_3B = INIT_3B;
defparam ram_inst.INIT_3C = INIT_3C;
defparam ram_inst.INIT_3D = INIT_3D;
defparam ram_inst.INIT_3E = INIT_3E;
defparam ram_inst.INIT_3F = INIT_3F;

`ifdef TIMINGCHECK
specify
   (RCLK *> RDATA[0]) = (1.0, 1.0);
   (RCLK *> RDATA[1]) = (1.0, 1.0);
   (RCLK *> RDATA[2]) = (1.0, 1.0);
   (RCLK *> RDATA[3]) = (1.0, 1.0);
   (RCLK *> RDATA[4]) = (1.0, 1.0);
   (RCLK *> RDATA[5]) = (1.0, 1.0);
   (RCLK *> RDATA[6]) = (1.0, 1.0);
   (RCLK *> RDATA[7]) = (1.0, 1.0);
   (RCLK *> RDATA[8]) = (1.0, 1.0);
   (RCLK *> RDATA[9]) = (1.0, 1.0);
   (RCLK *> RDATA[10]) = (1.0, 1.0);
   (RCLK *> RDATA[11]) = (1.0, 1.0);
   (RCLK *> RDATA[12]) = (1.0, 1.0);
   (RCLK *> RDATA[13]) = (1.0, 1.0);
   (RCLK *> RDATA[14]) = (1.0, 1.0);
   (RCLK *> RDATA[15]) = (1.0, 1.0);
   $setup(posedge MASK[0], posedge WCLK, 1.0);
   $setup(negedge MASK[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[0], 1.0);
   $hold(posedge WCLK, negedge MASK[0], 1.0);
   $setup(posedge MASK[1], posedge WCLK, 1.0);
   $setup(negedge MASK[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[1], 1.0);
   $hold(posedge WCLK, negedge MASK[1], 1.0);
   $setup(posedge MASK[2], posedge WCLK, 1.0);
   $setup(negedge MASK[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[2], 1.0);
   $hold(posedge WCLK, negedge MASK[2], 1.0);
   $setup(posedge MASK[3], posedge WCLK, 1.0);
   $setup(negedge MASK[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[3], 1.0);
   $hold(posedge WCLK, negedge MASK[3], 1.0);
   $setup(posedge MASK[4], posedge WCLK, 1.0);
   $setup(negedge MASK[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[4], 1.0);
   $hold(posedge WCLK, negedge MASK[4], 1.0);
   $setup(posedge MASK[5], posedge WCLK, 1.0);
   $setup(negedge MASK[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[5], 1.0);
   $hold(posedge WCLK, negedge MASK[5], 1.0);
   $setup(posedge MASK[6], posedge WCLK, 1.0);
   $setup(negedge MASK[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[6], 1.0);
   $hold(posedge WCLK, negedge MASK[6], 1.0);
   $setup(posedge MASK[7], posedge WCLK, 1.0);
   $setup(negedge MASK[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[7], 1.0);
   $hold(posedge WCLK, negedge MASK[7], 1.0);
   $setup(posedge MASK[8], posedge WCLK, 1.0);
   $setup(negedge MASK[8], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[8], 1.0);
   $hold(posedge WCLK, negedge MASK[8], 1.0);
   $setup(posedge MASK[9], posedge WCLK, 1.0);
   $setup(negedge MASK[9], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[9], 1.0);
   $hold(posedge WCLK, negedge MASK[9], 1.0);
   $setup(posedge MASK[10], posedge WCLK, 1.0);
   $setup(negedge MASK[10], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[10], 1.0);
   $hold(posedge WCLK, negedge MASK[10], 1.0);
   $setup(posedge MASK[11], posedge WCLK, 1.0);
   $setup(negedge MASK[11], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[11], 1.0);
   $hold(posedge WCLK, negedge MASK[11], 1.0);
   $setup(posedge MASK[12], posedge WCLK, 1.0);
   $setup(negedge MASK[12], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[12], 1.0);
   $hold(posedge WCLK, negedge MASK[12], 1.0);
   $setup(posedge MASK[13], posedge WCLK, 1.0);
   $setup(negedge MASK[13], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[13], 1.0);
   $hold(posedge WCLK, negedge MASK[13], 1.0);
   $setup(posedge MASK[14], posedge WCLK, 1.0);
   $setup(negedge MASK[14], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[14], 1.0);
   $hold(posedge WCLK, negedge MASK[14], 1.0);
   $setup(posedge MASK[15], posedge WCLK, 1.0);
   $setup(negedge MASK[15], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[15], 1.0);
   $hold(posedge WCLK, negedge MASK[15], 1.0);
   $setup(posedge WADDR[0], posedge WCLK, 1.0);
   $setup(negedge WADDR[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[0], 1.0);
   $hold(posedge WCLK, negedge WADDR[0], 1.0);
   $setup(posedge WADDR[1], posedge WCLK, 1.0);
   $setup(negedge WADDR[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[1], 1.0);
   $hold(posedge WCLK, negedge WADDR[1], 1.0);
   $setup(posedge WADDR[2], posedge WCLK, 1.0);
   $setup(negedge WADDR[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[2], 1.0);
   $hold(posedge WCLK, negedge WADDR[2], 1.0);
   $setup(posedge WADDR[3], posedge WCLK, 1.0);
   $setup(negedge WADDR[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[3], 1.0);
   $hold(posedge WCLK, negedge WADDR[3], 1.0);
   $setup(posedge WADDR[4], posedge WCLK, 1.0);
   $setup(negedge WADDR[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[4], 1.0);
   $hold(posedge WCLK, negedge WADDR[4], 1.0);
   $setup(posedge WADDR[5], posedge WCLK, 1.0);
   $setup(negedge WADDR[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[5], 1.0);
   $hold(posedge WCLK, negedge WADDR[5], 1.0);
   $setup(posedge WADDR[6], posedge WCLK, 1.0);
   $setup(negedge WADDR[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[6], 1.0);
   $hold(posedge WCLK, negedge WADDR[6], 1.0);
   $setup(posedge WADDR[7], posedge WCLK, 1.0);
   $setup(negedge WADDR[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[7], 1.0);
   $hold(posedge WCLK, negedge WADDR[7], 1.0);
   $setup(posedge WADDR[8], posedge WCLK, 1.0);
   $setup(negedge WADDR[8], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[8], 1.0);
   $hold(posedge WCLK, negedge WADDR[8], 1.0);
   $setup(posedge WADDR[9], posedge WCLK, 1.0);
   $setup(negedge WADDR[9], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[9], 1.0);
   $hold(posedge WCLK, negedge WADDR[9], 1.0);
   $setup(posedge WADDR[10], posedge WCLK, 1.0);
   $setup(negedge WADDR[10], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[10], 1.0);
   $hold(posedge WCLK, negedge WADDR[10], 1.0);
   $setup(posedge WADDR[11], posedge WCLK, 1.0);
   $setup(negedge WADDR[11], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[11], 1.0);
   $hold(posedge WCLK, negedge WADDR[11], 1.0);
   $setup(posedge WADDR[12], posedge WCLK, 1.0);
   $setup(negedge WADDR[12], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[12], 1.0);
   $hold(posedge WCLK, negedge WADDR[12], 1.0);
   $setup(posedge WDATA[0], posedge WCLK, 1.0);
   $setup(negedge WDATA[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[0], 1.0);
   $hold(posedge WCLK, negedge WDATA[0], 1.0);
   $setup(posedge WDATA[1], posedge WCLK, 1.0);
   $setup(negedge WDATA[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[1], 1.0);
   $hold(posedge WCLK, negedge WDATA[1], 1.0);
   $setup(posedge WDATA[2], posedge WCLK, 1.0);
   $setup(negedge WDATA[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[2], 1.0);
   $hold(posedge WCLK, negedge WDATA[2], 1.0);
   $setup(posedge WDATA[3], posedge WCLK, 1.0);
   $setup(negedge WDATA[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[3], 1.0);
   $hold(posedge WCLK, negedge WDATA[3], 1.0);
   $setup(posedge WDATA[4], posedge WCLK, 1.0);
   $setup(negedge WDATA[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[4], 1.0);
   $hold(posedge WCLK, negedge WDATA[4], 1.0);
   $setup(posedge WDATA[5], posedge WCLK, 1.0);
   $setup(negedge WDATA[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[5], 1.0);
   $hold(posedge WCLK, negedge WDATA[5], 1.0);
   $setup(posedge WDATA[6], posedge WCLK, 1.0);
   $setup(negedge WDATA[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[6], 1.0);
   $hold(posedge WCLK, negedge WDATA[6], 1.0);
   $setup(posedge WDATA[7], posedge WCLK, 1.0);
   $setup(negedge WDATA[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[7], 1.0);
   $hold(posedge WCLK, negedge WDATA[7], 1.0);
   $setup(posedge WDATA[8], posedge WCLK, 1.0);
   $setup(negedge WDATA[8], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[8], 1.0);
   $hold(posedge WCLK, negedge WDATA[8], 1.0);
   $setup(posedge WDATA[9], posedge WCLK, 1.0);
   $setup(negedge WDATA[9], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[9], 1.0);
   $hold(posedge WCLK, negedge WDATA[9], 1.0);
   $setup(posedge WDATA[10], posedge WCLK, 1.0);
   $setup(negedge WDATA[10], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[10], 1.0);
   $hold(posedge WCLK, negedge WDATA[10], 1.0);
   $setup(posedge WDATA[11], posedge WCLK, 1.0);
   $setup(negedge WDATA[11], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[11], 1.0);
   $hold(posedge WCLK, negedge WDATA[11], 1.0);
   $setup(posedge WDATA[12], posedge WCLK, 1.0);
   $setup(negedge WDATA[12], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[12], 1.0);
   $hold(posedge WCLK, negedge WDATA[12], 1.0);
   $setup(posedge WDATA[13], posedge WCLK, 1.0);
   $setup(negedge WDATA[13], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[13], 1.0);
   $hold(posedge WCLK, negedge WDATA[13], 1.0);
   $setup(posedge WDATA[14], posedge WCLK, 1.0);
   $setup(negedge WDATA[14], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[14], 1.0);
   $hold(posedge WCLK, negedge WDATA[14], 1.0);
   $setup(posedge WDATA[15], posedge WCLK, 1.0);
   $setup(negedge WDATA[15], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[15], 1.0);
   $hold(posedge WCLK, negedge WDATA[15], 1.0);
   $setup(posedge WCLKE, posedge WCLK, 1.0);
   $setup(negedge WCLKE, posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WCLKE, 1.0);
   $hold(posedge WCLK, negedge WCLKE, 1.0);
   $setup(posedge WE, posedge WCLK, 1.0);
   $setup(negedge WE, posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WE, 1.0);
   $hold(posedge WCLK, negedge WE, 1.0);
   $setup(posedge RADDR[0], posedge RCLK, 1.0);
   $setup(negedge RADDR[0], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[0], 1.0);
   $hold(posedge RCLK, negedge RADDR[0], 1.0);
   $setup(posedge RADDR[1], posedge RCLK, 1.0);
   $setup(negedge RADDR[1], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[1], 1.0);
   $hold(posedge RCLK, negedge RADDR[1], 1.0);
   $setup(posedge RADDR[2], posedge RCLK, 1.0);
   $setup(negedge RADDR[2], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[2], 1.0);
   $hold(posedge RCLK, negedge RADDR[2], 1.0);
   $setup(posedge RADDR[3], posedge RCLK, 1.0);
   $setup(negedge RADDR[3], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[3], 1.0);
   $hold(posedge RCLK, negedge RADDR[3], 1.0);
   $setup(posedge RADDR[4], posedge RCLK, 1.0);
   $setup(negedge RADDR[4], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[4], 1.0);
   $hold(posedge RCLK, negedge RADDR[4], 1.0);
   $setup(posedge RADDR[5], posedge RCLK, 1.0);
   $setup(negedge RADDR[5], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[5], 1.0);
   $hold(posedge RCLK, negedge RADDR[5], 1.0);
   $setup(posedge RADDR[6], posedge RCLK, 1.0);
   $setup(negedge RADDR[6], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[6], 1.0);
   $hold(posedge RCLK, negedge RADDR[6], 1.0);
   $setup(posedge RADDR[7], posedge RCLK, 1.0);
   $setup(negedge RADDR[7], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[7], 1.0);
   $hold(posedge RCLK, negedge RADDR[7], 1.0);
   $setup(posedge RADDR[8], posedge RCLK, 1.0);
   $setup(negedge RADDR[8], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[8], 1.0);
   $hold(posedge RCLK, negedge RADDR[8], 1.0);
   $setup(posedge RADDR[9], posedge RCLK, 1.0);
   $setup(negedge RADDR[9], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[9], 1.0);
   $hold(posedge RCLK, negedge RADDR[9], 1.0);
   $setup(posedge RADDR[10], posedge RCLK, 1.0);
   $setup(negedge RADDR[10], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[10], 1.0);
   $hold(posedge RCLK, negedge RADDR[10], 1.0);
   $setup(posedge RADDR[11], posedge RCLK, 1.0);
   $setup(negedge RADDR[11], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[11], 1.0);
   $hold(posedge RCLK, negedge RADDR[11], 1.0);
   $setup(posedge RADDR[12], posedge RCLK, 1.0);
   $setup(negedge RADDR[12], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[12], 1.0);
   $hold(posedge RCLK, negedge RADDR[12], 1.0);
   $setup(posedge RCLKE, posedge RCLK, 1.0);
   $setup(negedge RCLKE, posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RCLKE, 1.0);
   $hold(posedge RCLK, negedge RCLKE, 1.0);
   $setup(posedge RE, posedge RCLK, 1.0);
   $setup(negedge RE, posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RE, 1.0);
   $hold(posedge RCLK, negedge RE, 1.0);
endspecify
`endif

endmodule // SB_RAM40_16K;

//---------------------------------------
//	--- SB_RAM40_16KNR
//---------------------------------------

`timescale 1ps/1ps
module SB_RAM40_16KNR ( RDATA, RCLKN, RCLKE, RE, RADDR, WCLK, WCLKE, WE, WADDR, MASK, WDATA ); 

output	[15:0]	RDATA;  
input         	RCLKN;   
input           RCLKE; 
input           RE; 
input	[12:0]  RADDR; 
input           WCLK; 
input           WCLKE; 
input           WE; 
input 	[12:0]  WADDR; 
input 	[15:0]  MASK; 
input 	[15:0]	WDATA; 

parameter WRITE_MODE = 0;    // Configure Write Port as 1024x16 (0)/ 20148x8 (1)/ 4096x4 (2)/ 8192x2 (3)     
parameter READ_MODE  = 0;    // Configure Read  Port as 1024x16 (0)/ 20148x8 (1)/ 4096x4 (2)/ 8192x2 (3)

parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;


wire RCLK;
assign (weak0, weak1) RCLKE =1'b1 ;
assign (weak0, weak1) RE =1'b0 ;
assign (weak0, weak1) WCLKE =1'b1 ;
assign (weak0, weak1) WE =1'b0 ;
assign RCLK = ~RCLKN;

SB_RAM40_16K ram40mh_16K_nr_inst (
	.RDATA(RDATA),
	.RCLK(RCLK),
	.RCLKE(RCLKE),
	.RE(RE),
	.RADDR(RADDR),
	.WCLK(WCLK),
	.WCLKE(WCLKE),
	.WE(WE),
	.WADDR(WADDR),
	.MASK(MASK),
	.WDATA(WDATA));

defparam ram40mh_16K_nr_inst.WRITE_MODE = WRITE_MODE;
defparam ram40mh_16K_nr_inst.READ_MODE = READ_MODE;

defparam ram40mh_16K_nr_inst.INIT_0 = INIT_0;
defparam ram40mh_16K_nr_inst.INIT_1 = INIT_1;
defparam ram40mh_16K_nr_inst.INIT_2 = INIT_2;
defparam ram40mh_16K_nr_inst.INIT_3 = INIT_3;
defparam ram40mh_16K_nr_inst.INIT_4 = INIT_4;
defparam ram40mh_16K_nr_inst.INIT_5 = INIT_5;
defparam ram40mh_16K_nr_inst.INIT_6 = INIT_6;
defparam ram40mh_16K_nr_inst.INIT_7 = INIT_7;
defparam ram40mh_16K_nr_inst.INIT_8 = INIT_8;
defparam ram40mh_16K_nr_inst.INIT_9 = INIT_9;
defparam ram40mh_16K_nr_inst.INIT_A = INIT_A;
defparam ram40mh_16K_nr_inst.INIT_B = INIT_B;
defparam ram40mh_16K_nr_inst.INIT_C = INIT_C;
defparam ram40mh_16K_nr_inst.INIT_D = INIT_D;
defparam ram40mh_16K_nr_inst.INIT_E = INIT_E;
defparam ram40mh_16K_nr_inst.INIT_F = INIT_F;

defparam ram40mh_16K_nr_inst.INIT_0 = INIT_0;
defparam ram40mh_16K_nr_inst.INIT_1 = INIT_1;
defparam ram40mh_16K_nr_inst.INIT_2 = INIT_2;
defparam ram40mh_16K_nr_inst.INIT_3 = INIT_3;
defparam ram40mh_16K_nr_inst.INIT_4 = INIT_4;
defparam ram40mh_16K_nr_inst.INIT_5 = INIT_5;
defparam ram40mh_16K_nr_inst.INIT_6 = INIT_6;
defparam ram40mh_16K_nr_inst.INIT_7 = INIT_7;
defparam ram40mh_16K_nr_inst.INIT_8 = INIT_8;
defparam ram40mh_16K_nr_inst.INIT_9 = INIT_9;
defparam ram40mh_16K_nr_inst.INIT_A = INIT_A;
defparam ram40mh_16K_nr_inst.INIT_B = INIT_B;
defparam ram40mh_16K_nr_inst.INIT_C = INIT_C;
defparam ram40mh_16K_nr_inst.INIT_D = INIT_D;
defparam ram40mh_16K_nr_inst.INIT_E = INIT_E;
defparam ram40mh_16K_nr_inst.INIT_F = INIT_F;

defparam ram40mh_16K_nr_inst.INIT_0 = INIT_0;
defparam ram40mh_16K_nr_inst.INIT_1 = INIT_1;
defparam ram40mh_16K_nr_inst.INIT_2 = INIT_2;
defparam ram40mh_16K_nr_inst.INIT_3 = INIT_3;
defparam ram40mh_16K_nr_inst.INIT_4 = INIT_4;
defparam ram40mh_16K_nr_inst.INIT_5 = INIT_5;
defparam ram40mh_16K_nr_inst.INIT_6 = INIT_6;
defparam ram40mh_16K_nr_inst.INIT_7 = INIT_7;
defparam ram40mh_16K_nr_inst.INIT_8 = INIT_8;
defparam ram40mh_16K_nr_inst.INIT_9 = INIT_9;
defparam ram40mh_16K_nr_inst.INIT_A = INIT_A;
defparam ram40mh_16K_nr_inst.INIT_B = INIT_B;
defparam ram40mh_16K_nr_inst.INIT_C = INIT_C;
defparam ram40mh_16K_nr_inst.INIT_D = INIT_D;
defparam ram40mh_16K_nr_inst.INIT_E = INIT_E;
defparam ram40mh_16K_nr_inst.INIT_F = INIT_F;

defparam ram40mh_16K_nr_inst.INIT_0 = INIT_0;
defparam ram40mh_16K_nr_inst.INIT_1 = INIT_1;
defparam ram40mh_16K_nr_inst.INIT_2 = INIT_2;
defparam ram40mh_16K_nr_inst.INIT_3 = INIT_3;
defparam ram40mh_16K_nr_inst.INIT_4 = INIT_4;
defparam ram40mh_16K_nr_inst.INIT_5 = INIT_5;
defparam ram40mh_16K_nr_inst.INIT_6 = INIT_6;
defparam ram40mh_16K_nr_inst.INIT_7 = INIT_7;
defparam ram40mh_16K_nr_inst.INIT_8 = INIT_8;
defparam ram40mh_16K_nr_inst.INIT_9 = INIT_9;
defparam ram40mh_16K_nr_inst.INIT_A = INIT_A;
defparam ram40mh_16K_nr_inst.INIT_B = INIT_B;
defparam ram40mh_16K_nr_inst.INIT_C = INIT_C;
defparam ram40mh_16K_nr_inst.INIT_D = INIT_D;
defparam ram40mh_16K_nr_inst.INIT_E = INIT_E;
defparam ram40mh_16K_nr_inst.INIT_F = INIT_F;

`ifdef TIMINGCHECK
specify
   (RCLKN *> RDATA[0]) = (1.0, 1.0);
   (RCLKN *> RDATA[1]) = (1.0, 1.0);
   (RCLKN *> RDATA[2]) = (1.0, 1.0);
   (RCLKN *> RDATA[3]) = (1.0, 1.0);
   (RCLKN *> RDATA[4]) = (1.0, 1.0);
   (RCLKN *> RDATA[5]) = (1.0, 1.0);
   (RCLKN *> RDATA[6]) = (1.0, 1.0);
   (RCLKN *> RDATA[7]) = (1.0, 1.0);
   (RCLKN *> RDATA[8]) = (1.0, 1.0);
   (RCLKN *> RDATA[9]) = (1.0, 1.0);
   (RCLKN *> RDATA[10]) = (1.0, 1.0);
   (RCLKN *> RDATA[11]) = (1.0, 1.0);
   (RCLKN *> RDATA[12]) = (1.0, 1.0);
   (RCLKN *> RDATA[13]) = (1.0, 1.0);
   (RCLKN *> RDATA[14]) = (1.0, 1.0);
   (RCLKN *> RDATA[15]) = (1.0, 1.0);
   $setup(posedge MASK[0], posedge WCLK, 1.0);
   $setup(negedge MASK[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[0], 1.0);
   $hold(posedge WCLK, negedge MASK[0], 1.0);
   $setup(posedge MASK[1], posedge WCLK, 1.0);
   $setup(negedge MASK[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[1], 1.0);
   $hold(posedge WCLK, negedge MASK[1], 1.0);
   $setup(posedge MASK[2], posedge WCLK, 1.0);
   $setup(negedge MASK[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[2], 1.0);
   $hold(posedge WCLK, negedge MASK[2], 1.0);
   $setup(posedge MASK[3], posedge WCLK, 1.0);
   $setup(negedge MASK[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[3], 1.0);
   $hold(posedge WCLK, negedge MASK[3], 1.0);
   $setup(posedge MASK[4], posedge WCLK, 1.0);
   $setup(negedge MASK[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[4], 1.0);
   $hold(posedge WCLK, negedge MASK[4], 1.0);
   $setup(posedge MASK[5], posedge WCLK, 1.0);
   $setup(negedge MASK[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[5], 1.0);
   $hold(posedge WCLK, negedge MASK[5], 1.0);
   $setup(posedge MASK[6], posedge WCLK, 1.0);
   $setup(negedge MASK[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[6], 1.0);
   $hold(posedge WCLK, negedge MASK[6], 1.0);
   $setup(posedge MASK[7], posedge WCLK, 1.0);
   $setup(negedge MASK[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[7], 1.0);
   $hold(posedge WCLK, negedge MASK[7], 1.0);
   $setup(posedge MASK[8], posedge WCLK, 1.0);
   $setup(negedge MASK[8], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[8], 1.0);
   $hold(posedge WCLK, negedge MASK[8], 1.0);
   $setup(posedge MASK[9], posedge WCLK, 1.0);
   $setup(negedge MASK[9], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[9], 1.0);
   $hold(posedge WCLK, negedge MASK[9], 1.0);
   $setup(posedge MASK[10], posedge WCLK, 1.0);
   $setup(negedge MASK[10], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[10], 1.0);
   $hold(posedge WCLK, negedge MASK[10], 1.0);
   $setup(posedge MASK[11], posedge WCLK, 1.0);
   $setup(negedge MASK[11], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[11], 1.0);
   $hold(posedge WCLK, negedge MASK[11], 1.0);
   $setup(posedge MASK[12], posedge WCLK, 1.0);
   $setup(negedge MASK[12], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[12], 1.0);
   $hold(posedge WCLK, negedge MASK[12], 1.0);
   $setup(posedge MASK[13], posedge WCLK, 1.0);
   $setup(negedge MASK[13], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[13], 1.0);
   $hold(posedge WCLK, negedge MASK[13], 1.0);
   $setup(posedge MASK[14], posedge WCLK, 1.0);
   $setup(negedge MASK[14], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[14], 1.0);
   $hold(posedge WCLK, negedge MASK[14], 1.0);
   $setup(posedge MASK[15], posedge WCLK, 1.0);
   $setup(negedge MASK[15], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge MASK[15], 1.0);
   $hold(posedge WCLK, negedge MASK[15], 1.0);
   $setup(posedge WADDR[0], posedge WCLK, 1.0);
   $setup(negedge WADDR[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[0], 1.0);
   $hold(posedge WCLK, negedge WADDR[0], 1.0);
   $setup(posedge WADDR[1], posedge WCLK, 1.0);
   $setup(negedge WADDR[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[1], 1.0);
   $hold(posedge WCLK, negedge WADDR[1], 1.0);
   $setup(posedge WADDR[2], posedge WCLK, 1.0);
   $setup(negedge WADDR[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[2], 1.0);
   $hold(posedge WCLK, negedge WADDR[2], 1.0);
   $setup(posedge WADDR[3], posedge WCLK, 1.0);
   $setup(negedge WADDR[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[3], 1.0);
   $hold(posedge WCLK, negedge WADDR[3], 1.0);
   $setup(posedge WADDR[4], posedge WCLK, 1.0);
   $setup(negedge WADDR[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[4], 1.0);
   $hold(posedge WCLK, negedge WADDR[4], 1.0);
   $setup(posedge WADDR[5], posedge WCLK, 1.0);
   $setup(negedge WADDR[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[5], 1.0);
   $hold(posedge WCLK, negedge WADDR[5], 1.0);
   $setup(posedge WADDR[6], posedge WCLK, 1.0);
   $setup(negedge WADDR[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[6], 1.0);
   $hold(posedge WCLK, negedge WADDR[6], 1.0);
   $setup(posedge WADDR[7], posedge WCLK, 1.0);
   $setup(negedge WADDR[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[7], 1.0);
   $hold(posedge WCLK, negedge WADDR[7], 1.0);
   $setup(posedge WADDR[8], posedge WCLK, 1.0);
   $setup(negedge WADDR[8], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[8], 1.0);
   $hold(posedge WCLK, negedge WADDR[8], 1.0);
   $setup(posedge WADDR[9], posedge WCLK, 1.0);
   $setup(negedge WADDR[9], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[9], 1.0);
   $hold(posedge WCLK, negedge WADDR[9], 1.0);
   $setup(posedge WADDR[10], posedge WCLK, 1.0);
   $setup(negedge WADDR[10], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[10], 1.0);
   $hold(posedge WCLK, negedge WADDR[10], 1.0);
   $setup(posedge WADDR[11], posedge WCLK, 1.0);
   $setup(negedge WADDR[11], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[11], 1.0);
   $hold(posedge WCLK, negedge WADDR[11], 1.0);
   $setup(posedge WADDR[12], posedge WCLK, 1.0);
   $setup(negedge WADDR[12], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WADDR[12], 1.0);
   $hold(posedge WCLK, negedge WADDR[12], 1.0);
   $setup(posedge WDATA[0], posedge WCLK, 1.0);
   $setup(negedge WDATA[0], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[0], 1.0);
   $hold(posedge WCLK, negedge WDATA[0], 1.0);
   $setup(posedge WDATA[1], posedge WCLK, 1.0);
   $setup(negedge WDATA[1], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[1], 1.0);
   $hold(posedge WCLK, negedge WDATA[1], 1.0);
   $setup(posedge WDATA[2], posedge WCLK, 1.0);
   $setup(negedge WDATA[2], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[2], 1.0);
   $hold(posedge WCLK, negedge WDATA[2], 1.0);
   $setup(posedge WDATA[3], posedge WCLK, 1.0);
   $setup(negedge WDATA[3], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[3], 1.0);
   $hold(posedge WCLK, negedge WDATA[3], 1.0);
   $setup(posedge WDATA[4], posedge WCLK, 1.0);
   $setup(negedge WDATA[4], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[4], 1.0);
   $hold(posedge WCLK, negedge WDATA[4], 1.0);
   $setup(posedge WDATA[5], posedge WCLK, 1.0);
   $setup(negedge WDATA[5], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[5], 1.0);
   $hold(posedge WCLK, negedge WDATA[5], 1.0);
   $setup(posedge WDATA[6], posedge WCLK, 1.0);
   $setup(negedge WDATA[6], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[6], 1.0);
   $hold(posedge WCLK, negedge WDATA[6], 1.0);
   $setup(posedge WDATA[7], posedge WCLK, 1.0);
   $setup(negedge WDATA[7], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[7], 1.0);
   $hold(posedge WCLK, negedge WDATA[7], 1.0);
   $setup(posedge WDATA[8], posedge WCLK, 1.0);
   $setup(negedge WDATA[8], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[8], 1.0);
   $hold(posedge WCLK, negedge WDATA[8], 1.0);
   $setup(posedge WDATA[9], posedge WCLK, 1.0);
   $setup(negedge WDATA[9], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[9], 1.0);
   $hold(posedge WCLK, negedge WDATA[9], 1.0);
   $setup(posedge WDATA[10], posedge WCLK, 1.0);
   $setup(negedge WDATA[10], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[10], 1.0);
   $hold(posedge WCLK, negedge WDATA[10], 1.0);
   $setup(posedge WDATA[11], posedge WCLK, 1.0);
   $setup(negedge WDATA[11], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[11], 1.0);
   $hold(posedge WCLK, negedge WDATA[11], 1.0);
   $setup(posedge WDATA[12], posedge WCLK, 1.0);
   $setup(negedge WDATA[12], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[12], 1.0);
   $hold(posedge WCLK, negedge WDATA[12], 1.0);
   $setup(posedge WDATA[13], posedge WCLK, 1.0);
   $setup(negedge WDATA[13], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[13], 1.0);
   $hold(posedge WCLK, negedge WDATA[13], 1.0);
   $setup(posedge WDATA[14], posedge WCLK, 1.0);
   $setup(negedge WDATA[14], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[14], 1.0);
   $hold(posedge WCLK, negedge WDATA[14], 1.0);
   $setup(posedge WDATA[15], posedge WCLK, 1.0);
   $setup(negedge WDATA[15], posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WDATA[15], 1.0);
   $hold(posedge WCLK, negedge WDATA[15], 1.0);
   $setup(posedge WCLKE, posedge WCLK, 1.0);
   $setup(negedge WCLKE, posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WCLKE, 1.0);
   $hold(posedge WCLK, negedge WCLKE, 1.0);
   $setup(posedge WE, posedge WCLK, 1.0);
   $setup(negedge WE, posedge WCLK, 1.0);
   $hold(posedge WCLK, posedge WE, 1.0);
   $hold(posedge WCLK, negedge WE, 1.0);
   $setup(posedge RADDR[0], posedge RCLKN, 1.0);
   $setup(negedge RADDR[0], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[0], 1.0);
   $hold(posedge RCLKN, negedge RADDR[0], 1.0);
   $setup(posedge RADDR[1], posedge RCLKN, 1.0);
   $setup(negedge RADDR[1], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[1], 1.0);
   $hold(posedge RCLKN, negedge RADDR[1], 1.0);
   $setup(posedge RADDR[2], posedge RCLKN, 1.0);
   $setup(negedge RADDR[2], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[2], 1.0);
   $hold(posedge RCLKN, negedge RADDR[2], 1.0);
   $setup(posedge RADDR[3], posedge RCLKN, 1.0);
   $setup(negedge RADDR[3], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[3], 1.0);
   $hold(posedge RCLKN, negedge RADDR[3], 1.0);
   $setup(posedge RADDR[4], posedge RCLKN, 1.0);
   $setup(negedge RADDR[4], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[4], 1.0);
   $hold(posedge RCLKN, negedge RADDR[4], 1.0);
   $setup(posedge RADDR[5], posedge RCLKN, 1.0);
   $setup(negedge RADDR[5], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[5], 1.0);
   $hold(posedge RCLKN, negedge RADDR[5], 1.0);
   $setup(posedge RADDR[6], posedge RCLKN, 1.0);
   $setup(negedge RADDR[6], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[6], 1.0);
   $hold(posedge RCLKN, negedge RADDR[6], 1.0);
   $setup(posedge RADDR[7], posedge RCLKN, 1.0);
   $setup(negedge RADDR[7], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[7], 1.0);
   $hold(posedge RCLKN, negedge RADDR[7], 1.0);
   $setup(posedge RADDR[8], posedge RCLKN, 1.0);
   $setup(negedge RADDR[8], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[8], 1.0);
   $hold(posedge RCLKN, negedge RADDR[8], 1.0);
   $setup(posedge RADDR[9], posedge RCLKN, 1.0);
   $setup(negedge RADDR[9], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[9], 1.0);
   $hold(posedge RCLKN, negedge RADDR[9], 1.0);
   $setup(posedge RADDR[10], posedge RCLKN, 1.0);
   $setup(negedge RADDR[10], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[10], 1.0);
   $hold(posedge RCLKN, negedge RADDR[10], 1.0);
   $setup(posedge RADDR[11], posedge RCLKN, 1.0);
   $setup(negedge RADDR[11], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[11], 1.0);
   $hold(posedge RCLKN, negedge RADDR[11], 1.0);
   $setup(posedge RADDR[12], posedge RCLKN, 1.0);
   $setup(negedge RADDR[12], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[12], 1.0);
   $hold(posedge RCLKN, negedge RADDR[12], 1.0);
   $setup(posedge RCLKE, posedge RCLKN, 1.0);
   $setup(negedge RCLKE, posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RCLKE, 1.0);
   $hold(posedge RCLKN, negedge RCLKE, 1.0);
   $setup(posedge RE, posedge RCLKN, 1.0);
   $setup(negedge RE, posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RE, 1.0);
   $hold(posedge RCLKN, negedge RE, 1.0);
endspecify
`endif
 
endmodule  // SB_RAM40_16KNR 

//---------------------------------------
//	--- SB_RAM40_16KNW
//---------------------------------------
`timescale 1ps/1ps
module  SB_RAM40_16KNW ( RDATA, RCLK, RCLKE, RE, RADDR, WCLKN, WCLKE, WE, WADDR, MASK, WDATA ); 

output	[15:0]	RDATA;  
input         	RCLK;   
input           RCLKE; 
input           RE; 
input	[12:0]  RADDR; 
input           WCLKN; 
input           WCLKE; 
input           WE; 
input 	[12:0]  WADDR; 
input 	[15:0]  MASK; 
input 	[15:0]	WDATA; 

parameter WRITE_MODE = 0;    // Configure Write Port as 1024x16 (0)/ 20148x8 (1)/ 4096x4 (2)/ 8192x2 (3)     
parameter READ_MODE  = 0;    // Configure Read  Port as 1024x16 (0)/ 20148x8 (1)/ 4096x4 (2)/ 8192x2 (3)

parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;


wire WCLK;
assign (weak0, weak1) RCLKE =1'b1 ;
assign (weak0, weak1) RE =1'b0 ;
assign (weak0, weak1) WCLKE =1'b1 ;
assign (weak0, weak1) WE =1'b0 ;
assign WCLK = ~WCLKN;

SB_RAM40_16K ram40mh_16K_nw_inst (
	.RDATA(RDATA),
	.RCLK(RCLK),
	.RCLKE(RCLKE),
	.RE(RE),
	.RADDR(RADDR),
	.WCLK(WCLK),
	.WCLKE(WCLKE),
	.WE(WE),
	.WADDR(WADDR),
	.MASK(MASK),
	.WDATA(WDATA));

defparam ram40mh_16K_nw_inst.WRITE_MODE = WRITE_MODE;
defparam ram40mh_16K_nw_inst.READ_MODE = READ_MODE;

defparam ram40mh_16K_nw_inst.INIT_0 = INIT_0;
defparam ram40mh_16K_nw_inst.INIT_1 = INIT_1;
defparam ram40mh_16K_nw_inst.INIT_2 = INIT_2;
defparam ram40mh_16K_nw_inst.INIT_3 = INIT_3;
defparam ram40mh_16K_nw_inst.INIT_4 = INIT_4;
defparam ram40mh_16K_nw_inst.INIT_5 = INIT_5;
defparam ram40mh_16K_nw_inst.INIT_6 = INIT_6;
defparam ram40mh_16K_nw_inst.INIT_7 = INIT_7;
defparam ram40mh_16K_nw_inst.INIT_8 = INIT_8;
defparam ram40mh_16K_nw_inst.INIT_9 = INIT_9;
defparam ram40mh_16K_nw_inst.INIT_A = INIT_A;
defparam ram40mh_16K_nw_inst.INIT_B = INIT_B;
defparam ram40mh_16K_nw_inst.INIT_C = INIT_C;
defparam ram40mh_16K_nw_inst.INIT_D = INIT_D;
defparam ram40mh_16K_nw_inst.INIT_E = INIT_E;
defparam ram40mh_16K_nw_inst.INIT_F = INIT_F;

defparam ram40mh_16K_nw_inst.INIT_0 = INIT_0;
defparam ram40mh_16K_nw_inst.INIT_1 = INIT_1;
defparam ram40mh_16K_nw_inst.INIT_2 = INIT_2;
defparam ram40mh_16K_nw_inst.INIT_3 = INIT_3;
defparam ram40mh_16K_nw_inst.INIT_4 = INIT_4;
defparam ram40mh_16K_nw_inst.INIT_5 = INIT_5;
defparam ram40mh_16K_nw_inst.INIT_6 = INIT_6;
defparam ram40mh_16K_nw_inst.INIT_7 = INIT_7;
defparam ram40mh_16K_nw_inst.INIT_8 = INIT_8;
defparam ram40mh_16K_nw_inst.INIT_9 = INIT_9;
defparam ram40mh_16K_nw_inst.INIT_A = INIT_A;
defparam ram40mh_16K_nw_inst.INIT_B = INIT_B;
defparam ram40mh_16K_nw_inst.INIT_C = INIT_C;
defparam ram40mh_16K_nw_inst.INIT_D = INIT_D;
defparam ram40mh_16K_nw_inst.INIT_E = INIT_E;
defparam ram40mh_16K_nw_inst.INIT_F = INIT_F;

defparam ram40mh_16K_nw_inst.INIT_0 = INIT_0;
defparam ram40mh_16K_nw_inst.INIT_1 = INIT_1;
defparam ram40mh_16K_nw_inst.INIT_2 = INIT_2;
defparam ram40mh_16K_nw_inst.INIT_3 = INIT_3;
defparam ram40mh_16K_nw_inst.INIT_4 = INIT_4;
defparam ram40mh_16K_nw_inst.INIT_5 = INIT_5;
defparam ram40mh_16K_nw_inst.INIT_6 = INIT_6;
defparam ram40mh_16K_nw_inst.INIT_7 = INIT_7;
defparam ram40mh_16K_nw_inst.INIT_8 = INIT_8;
defparam ram40mh_16K_nw_inst.INIT_9 = INIT_9;
defparam ram40mh_16K_nw_inst.INIT_A = INIT_A;
defparam ram40mh_16K_nw_inst.INIT_B = INIT_B;
defparam ram40mh_16K_nw_inst.INIT_C = INIT_C;
defparam ram40mh_16K_nw_inst.INIT_D = INIT_D;
defparam ram40mh_16K_nw_inst.INIT_E = INIT_E;
defparam ram40mh_16K_nw_inst.INIT_F = INIT_F;

defparam ram40mh_16K_nw_inst.INIT_0 = INIT_0;
defparam ram40mh_16K_nw_inst.INIT_1 = INIT_1;
defparam ram40mh_16K_nw_inst.INIT_2 = INIT_2;
defparam ram40mh_16K_nw_inst.INIT_3 = INIT_3;
defparam ram40mh_16K_nw_inst.INIT_4 = INIT_4;
defparam ram40mh_16K_nw_inst.INIT_5 = INIT_5;
defparam ram40mh_16K_nw_inst.INIT_6 = INIT_6;
defparam ram40mh_16K_nw_inst.INIT_7 = INIT_7;
defparam ram40mh_16K_nw_inst.INIT_8 = INIT_8;
defparam ram40mh_16K_nw_inst.INIT_9 = INIT_9;
defparam ram40mh_16K_nw_inst.INIT_A = INIT_A;
defparam ram40mh_16K_nw_inst.INIT_B = INIT_B;
defparam ram40mh_16K_nw_inst.INIT_C = INIT_C;
defparam ram40mh_16K_nw_inst.INIT_D = INIT_D;
defparam ram40mh_16K_nw_inst.INIT_E = INIT_E;
defparam ram40mh_16K_nw_inst.INIT_F = INIT_F;

`ifdef TIMINGCHECK
specify
   (RCLK *> RDATA[0]) = (1.0, 1.0);
   (RCLK *> RDATA[1]) = (1.0, 1.0);
   (RCLK *> RDATA[2]) = (1.0, 1.0);
   (RCLK *> RDATA[3]) = (1.0, 1.0);
   (RCLK *> RDATA[4]) = (1.0, 1.0);
   (RCLK *> RDATA[5]) = (1.0, 1.0);
   (RCLK *> RDATA[6]) = (1.0, 1.0);
   (RCLK *> RDATA[7]) = (1.0, 1.0);
   (RCLK *> RDATA[8]) = (1.0, 1.0);
   (RCLK *> RDATA[9]) = (1.0, 1.0);
   (RCLK *> RDATA[10]) = (1.0, 1.0);
   (RCLK *> RDATA[11]) = (1.0, 1.0);
   (RCLK *> RDATA[12]) = (1.0, 1.0);
   (RCLK *> RDATA[13]) = (1.0, 1.0);
   (RCLK *> RDATA[14]) = (1.0, 1.0);
   (RCLK *> RDATA[15]) = (1.0, 1.0);
   $setup(posedge MASK[0], posedge WCLKN, 1.0);
   $setup(negedge MASK[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[0], 1.0);
   $hold(posedge WCLKN, negedge MASK[0], 1.0);
   $setup(posedge MASK[1], posedge WCLKN, 1.0);
   $setup(negedge MASK[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[1], 1.0);
   $hold(posedge WCLKN, negedge MASK[1], 1.0);
   $setup(posedge MASK[2], posedge WCLKN, 1.0);
   $setup(negedge MASK[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[2], 1.0);
   $hold(posedge WCLKN, negedge MASK[2], 1.0);
   $setup(posedge MASK[3], posedge WCLKN, 1.0);
   $setup(negedge MASK[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[3], 1.0);
   $hold(posedge WCLKN, negedge MASK[3], 1.0);
   $setup(posedge MASK[4], posedge WCLKN, 1.0);
   $setup(negedge MASK[4], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[4], 1.0);
   $hold(posedge WCLKN, negedge MASK[4], 1.0);
   $setup(posedge MASK[5], posedge WCLKN, 1.0);
   $setup(negedge MASK[5], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[5], 1.0);
   $hold(posedge WCLKN, negedge MASK[5], 1.0);
   $setup(posedge MASK[6], posedge WCLKN, 1.0);
   $setup(negedge MASK[6], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[6], 1.0);
   $hold(posedge WCLKN, negedge MASK[6], 1.0);
   $setup(posedge MASK[7], posedge WCLKN, 1.0);
   $setup(negedge MASK[7], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[7], 1.0);
   $hold(posedge WCLKN, negedge MASK[7], 1.0);
   $setup(posedge MASK[8], posedge WCLKN, 1.0);
   $setup(negedge MASK[8], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[8], 1.0);
   $hold(posedge WCLKN, negedge MASK[8], 1.0);
   $setup(posedge MASK[9], posedge WCLKN, 1.0);
   $setup(negedge MASK[9], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[9], 1.0);
   $hold(posedge WCLKN, negedge MASK[9], 1.0);
   $setup(posedge MASK[10], posedge WCLKN, 1.0);
   $setup(negedge MASK[10], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[10], 1.0);
   $hold(posedge WCLKN, negedge MASK[10], 1.0);
   $setup(posedge MASK[11], posedge WCLKN, 1.0);
   $setup(negedge MASK[11], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[11], 1.0);
   $hold(posedge WCLKN, negedge MASK[11], 1.0);
   $setup(posedge MASK[12], posedge WCLKN, 1.0);
   $setup(negedge MASK[12], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[12], 1.0);
   $hold(posedge WCLKN, negedge MASK[12], 1.0);
   $setup(posedge MASK[13], posedge WCLKN, 1.0);
   $setup(negedge MASK[13], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[13], 1.0);
   $hold(posedge WCLKN, negedge MASK[13], 1.0);
   $setup(posedge MASK[14], posedge WCLKN, 1.0);
   $setup(negedge MASK[14], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[14], 1.0);
   $hold(posedge WCLKN, negedge MASK[14], 1.0);
   $setup(posedge MASK[15], posedge WCLKN, 1.0);
   $setup(negedge MASK[15], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[15], 1.0);
   $hold(posedge WCLKN, negedge MASK[15], 1.0);
   $setup(posedge WADDR[0], posedge WCLKN, 1.0);
   $setup(negedge WADDR[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[0], 1.0);
   $hold(posedge WCLKN, negedge WADDR[0], 1.0);
   $setup(posedge WADDR[1], posedge WCLKN, 1.0);
   $setup(negedge WADDR[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[1], 1.0);
   $hold(posedge WCLKN, negedge WADDR[1], 1.0);
   $setup(posedge WADDR[2], posedge WCLKN, 1.0);
   $setup(negedge WADDR[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[2], 1.0);
   $hold(posedge WCLKN, negedge WADDR[2], 1.0);
   $setup(posedge WADDR[3], posedge WCLKN, 1.0);
   $setup(negedge WADDR[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[3], 1.0);
   $hold(posedge WCLKN, negedge WADDR[3], 1.0);
   $setup(posedge WADDR[4], posedge WCLKN, 1.0);
   $setup(negedge WADDR[4], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[4], 1.0);
   $hold(posedge WCLKN, negedge WADDR[4], 1.0);
   $setup(posedge WADDR[5], posedge WCLKN, 1.0);
   $setup(negedge WADDR[5], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[5], 1.0);
   $hold(posedge WCLKN, negedge WADDR[5], 1.0);
   $setup(posedge WADDR[6], posedge WCLKN, 1.0);
   $setup(negedge WADDR[6], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[6], 1.0);
   $hold(posedge WCLKN, negedge WADDR[6], 1.0);
   $setup(posedge WADDR[7], posedge WCLKN, 1.0);
   $setup(negedge WADDR[7], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[7], 1.0);
   $hold(posedge WCLKN, negedge WADDR[7], 1.0);
   $setup(posedge WADDR[8], posedge WCLKN, 1.0);
   $setup(negedge WADDR[8], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[8], 1.0);
   $hold(posedge WCLKN, negedge WADDR[8], 1.0);
   $setup(posedge WADDR[9], posedge WCLKN, 1.0);
   $setup(negedge WADDR[9], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[9], 1.0);
   $hold(posedge WCLKN, negedge WADDR[9], 1.0);
   $setup(posedge WADDR[10], posedge WCLKN, 1.0);
   $setup(negedge WADDR[10], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[10], 1.0);
   $hold(posedge WCLKN, negedge WADDR[10], 1.0);
   $setup(posedge WADDR[11], posedge WCLKN, 1.0);
   $setup(negedge WADDR[11], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[11], 1.0);
   $hold(posedge WCLKN, negedge WADDR[11], 1.0);
   $setup(posedge WADDR[12], posedge WCLKN, 1.0);
   $setup(negedge WADDR[12], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[12], 1.0);
   $hold(posedge WCLKN, negedge WADDR[12], 1.0);
   $setup(posedge WDATA[0], posedge WCLKN, 1.0);
   $setup(negedge WDATA[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[0], 1.0);
   $hold(posedge WCLKN, negedge WDATA[0], 1.0);
   $setup(posedge WDATA[1], posedge WCLKN, 1.0);
   $setup(negedge WDATA[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[1], 1.0);
   $hold(posedge WCLKN, negedge WDATA[1], 1.0);
   $setup(posedge WDATA[2], posedge WCLKN, 1.0);
   $setup(negedge WDATA[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[2], 1.0);
   $hold(posedge WCLKN, negedge WDATA[2], 1.0);
   $setup(posedge WDATA[3], posedge WCLKN, 1.0);
   $setup(negedge WDATA[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[3], 1.0);
   $hold(posedge WCLKN, negedge WDATA[3], 1.0);
   $setup(posedge WDATA[4], posedge WCLKN, 1.0);
   $setup(negedge WDATA[4], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[4], 1.0);
   $hold(posedge WCLKN, negedge WDATA[4], 1.0);
   $setup(posedge WDATA[5], posedge WCLKN, 1.0);
   $setup(negedge WDATA[5], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[5], 1.0);
   $hold(posedge WCLKN, negedge WDATA[5], 1.0);
   $setup(posedge WDATA[6], posedge WCLKN, 1.0);
   $setup(negedge WDATA[6], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[6], 1.0);
   $hold(posedge WCLKN, negedge WDATA[6], 1.0);
   $setup(posedge WDATA[7], posedge WCLKN, 1.0);
   $setup(negedge WDATA[7], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[7], 1.0);
   $hold(posedge WCLKN, negedge WDATA[7], 1.0);
   $setup(posedge WDATA[8], posedge WCLKN, 1.0);
   $setup(negedge WDATA[8], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[8], 1.0);
   $hold(posedge WCLKN, negedge WDATA[8], 1.0);
   $setup(posedge WDATA[9], posedge WCLKN, 1.0);
   $setup(negedge WDATA[9], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[9], 1.0);
   $hold(posedge WCLKN, negedge WDATA[9], 1.0);
   $setup(posedge WDATA[10], posedge WCLKN, 1.0);
   $setup(negedge WDATA[10], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[10], 1.0);
   $hold(posedge WCLKN, negedge WDATA[10], 1.0);
   $setup(posedge WDATA[11], posedge WCLKN, 1.0);
   $setup(negedge WDATA[11], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[11], 1.0);
   $hold(posedge WCLKN, negedge WDATA[11], 1.0);
   $setup(posedge WDATA[12], posedge WCLKN, 1.0);
   $setup(negedge WDATA[12], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[12], 1.0);
   $hold(posedge WCLKN, negedge WDATA[12], 1.0);
   $setup(posedge WDATA[13], posedge WCLKN, 1.0);
   $setup(negedge WDATA[13], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[13], 1.0);
   $hold(posedge WCLKN, negedge WDATA[13], 1.0);
   $setup(posedge WDATA[14], posedge WCLKN, 1.0);
   $setup(negedge WDATA[14], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[14], 1.0);
   $hold(posedge WCLKN, negedge WDATA[14], 1.0);
   $setup(posedge WDATA[15], posedge WCLKN, 1.0);
   $setup(negedge WDATA[15], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[15], 1.0);
   $hold(posedge WCLKN, negedge WDATA[15], 1.0);
   $setup(posedge WCLKE, posedge WCLKN, 1.0);
   $setup(negedge WCLKE, posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WCLKE, 1.0);
   $hold(posedge WCLKN, negedge WCLKE, 1.0);
   $setup(posedge WE, posedge WCLKN, 1.0);
   $setup(negedge WE, posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WE, 1.0);
   $hold(posedge WCLKN, negedge WE, 1.0);
   $setup(posedge RADDR[0], posedge RCLK, 1.0);
   $setup(negedge RADDR[0], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[0], 1.0);
   $hold(posedge RCLK, negedge RADDR[0], 1.0);
   $setup(posedge RADDR[1], posedge RCLK, 1.0);
   $setup(negedge RADDR[1], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[1], 1.0);
   $hold(posedge RCLK, negedge RADDR[1], 1.0);
   $setup(posedge RADDR[2], posedge RCLK, 1.0);
   $setup(negedge RADDR[2], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[2], 1.0);
   $hold(posedge RCLK, negedge RADDR[2], 1.0);
   $setup(posedge RADDR[3], posedge RCLK, 1.0);
   $setup(negedge RADDR[3], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[3], 1.0);
   $hold(posedge RCLK, negedge RADDR[3], 1.0);
   $setup(posedge RADDR[4], posedge RCLK, 1.0);
   $setup(negedge RADDR[4], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[4], 1.0);
   $hold(posedge RCLK, negedge RADDR[4], 1.0);
   $setup(posedge RADDR[5], posedge RCLK, 1.0);
   $setup(negedge RADDR[5], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[5], 1.0);
   $hold(posedge RCLK, negedge RADDR[5], 1.0);
   $setup(posedge RADDR[6], posedge RCLK, 1.0);
   $setup(negedge RADDR[6], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[6], 1.0);
   $hold(posedge RCLK, negedge RADDR[6], 1.0);
   $setup(posedge RADDR[7], posedge RCLK, 1.0);
   $setup(negedge RADDR[7], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[7], 1.0);
   $hold(posedge RCLK, negedge RADDR[7], 1.0);
   $setup(posedge RADDR[8], posedge RCLK, 1.0);
   $setup(negedge RADDR[8], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[8], 1.0);
   $hold(posedge RCLK, negedge RADDR[8], 1.0);
   $setup(posedge RADDR[9], posedge RCLK, 1.0);
   $setup(negedge RADDR[9], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[9], 1.0);
   $hold(posedge RCLK, negedge RADDR[9], 1.0);
   $setup(posedge RADDR[10], posedge RCLK, 1.0);
   $setup(negedge RADDR[10], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[10], 1.0);
   $hold(posedge RCLK, negedge RADDR[10], 1.0);
   $setup(posedge RADDR[11], posedge RCLK, 1.0);
   $setup(negedge RADDR[11], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[11], 1.0);
   $hold(posedge RCLK, negedge RADDR[11], 1.0);
   $setup(posedge RADDR[12], posedge RCLK, 1.0);
   $setup(negedge RADDR[12], posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RADDR[12], 1.0);
   $hold(posedge RCLK, negedge RADDR[12], 1.0);
   $setup(posedge RCLKE, posedge RCLK, 1.0);
   $setup(negedge RCLKE, posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RCLKE, 1.0);
   $hold(posedge RCLK, negedge RCLKE, 1.0);
   $setup(posedge RE, posedge RCLK, 1.0);
   $setup(negedge RE, posedge RCLK, 1.0);
   $hold(posedge RCLK, posedge RE, 1.0);
   $hold(posedge RCLK, negedge RE, 1.0);
endspecify
`endif
  
endmodule  // SB_RAM40_16KNW

// ---------------------------------------
// 	--- SB_RAM40_16KNRNW
// ---------------------------------------
`timescale 1ps/1ps
module SB_RAM40_16KNRNW ( RDATA, RCLKN, RCLKE, RE, RADDR, WCLKN, WCLKE, WE, WADDR, MASK, WDATA );  

output	[15:0]	RDATA;  
input         	RCLKN;   
input           RCLKE; 
input           RE; 
input	[12:0]  RADDR; 
input           WCLKN; 
input           WCLKE; 
input           WE; 
input 	[12:0]  WADDR; 
input 	[15:0]  MASK; 
input 	[15:0]	WDATA; 

parameter WRITE_MODE = 0;    // Configure Write Port as 1024x16 (0)/ 20148x8 (1)/ 4096x4 (2)/ 8192x2 (3)     
parameter READ_MODE  = 0;    // Configure Read  Port as 1024x16 (0)/ 20148x8 (1)/ 4096x4 (2)/ 8192x2 (3)

parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;   


wire RCLK;
wire WCLK; 
assign (weak0, weak1) RCLKE =1'b1 ;
assign (weak0, weak1) RE =1'b0 ;
assign (weak0, weak1) WCLKE =1'b1 ;
assign (weak0, weak1) WE =1'b0 ;
assign RCLK = ~RCLKN;
assign WCLK = ~WCLKN; 

SB_RAM40_16K ram40mh_16K_nrnw_inst (
	.RDATA(RDATA),
	.RCLK(RCLK),
	.RCLKE(RCLKE),
	.RE(RE),
	.RADDR(RADDR),
	.WCLK(WCLK),
	.WCLKE(WCLKE),
	.WE(WE),
	.WADDR(WADDR),
	.MASK(MASK),
	.WDATA(WDATA));

defparam ram40mh_16K_nrnw_inst.WRITE_MODE = WRITE_MODE;
defparam ram40mh_16K_nrnw_inst.READ_MODE = READ_MODE;

defparam ram40mh_16K_nrnw_inst.INIT_0 = INIT_0;
defparam ram40mh_16K_nrnw_inst.INIT_1 = INIT_1;
defparam ram40mh_16K_nrnw_inst.INIT_2 = INIT_2;
defparam ram40mh_16K_nrnw_inst.INIT_3 = INIT_3;
defparam ram40mh_16K_nrnw_inst.INIT_4 = INIT_4;
defparam ram40mh_16K_nrnw_inst.INIT_5 = INIT_5;
defparam ram40mh_16K_nrnw_inst.INIT_6 = INIT_6;
defparam ram40mh_16K_nrnw_inst.INIT_7 = INIT_7;
defparam ram40mh_16K_nrnw_inst.INIT_8 = INIT_8;
defparam ram40mh_16K_nrnw_inst.INIT_9 = INIT_9;
defparam ram40mh_16K_nrnw_inst.INIT_A = INIT_A;
defparam ram40mh_16K_nrnw_inst.INIT_B = INIT_B;
defparam ram40mh_16K_nrnw_inst.INIT_C = INIT_C;
defparam ram40mh_16K_nrnw_inst.INIT_D = INIT_D;
defparam ram40mh_16K_nrnw_inst.INIT_E = INIT_E;
defparam ram40mh_16K_nrnw_inst.INIT_F = INIT_F;

defparam ram40mh_16K_nrnw_inst.INIT_0 = INIT_0;
defparam ram40mh_16K_nrnw_inst.INIT_1 = INIT_1;
defparam ram40mh_16K_nrnw_inst.INIT_2 = INIT_2;
defparam ram40mh_16K_nrnw_inst.INIT_3 = INIT_3;
defparam ram40mh_16K_nrnw_inst.INIT_4 = INIT_4;
defparam ram40mh_16K_nrnw_inst.INIT_5 = INIT_5;
defparam ram40mh_16K_nrnw_inst.INIT_6 = INIT_6;
defparam ram40mh_16K_nrnw_inst.INIT_7 = INIT_7;
defparam ram40mh_16K_nrnw_inst.INIT_8 = INIT_8;
defparam ram40mh_16K_nrnw_inst.INIT_9 = INIT_9;
defparam ram40mh_16K_nrnw_inst.INIT_A = INIT_A;
defparam ram40mh_16K_nrnw_inst.INIT_B = INIT_B;
defparam ram40mh_16K_nrnw_inst.INIT_C = INIT_C;
defparam ram40mh_16K_nrnw_inst.INIT_D = INIT_D;
defparam ram40mh_16K_nrnw_inst.INIT_E = INIT_E;
defparam ram40mh_16K_nrnw_inst.INIT_F = INIT_F;

defparam ram40mh_16K_nrnw_inst.INIT_0 = INIT_0;
defparam ram40mh_16K_nrnw_inst.INIT_1 = INIT_1;
defparam ram40mh_16K_nrnw_inst.INIT_2 = INIT_2;
defparam ram40mh_16K_nrnw_inst.INIT_3 = INIT_3;
defparam ram40mh_16K_nrnw_inst.INIT_4 = INIT_4;
defparam ram40mh_16K_nrnw_inst.INIT_5 = INIT_5;
defparam ram40mh_16K_nrnw_inst.INIT_6 = INIT_6;
defparam ram40mh_16K_nrnw_inst.INIT_7 = INIT_7;
defparam ram40mh_16K_nrnw_inst.INIT_8 = INIT_8;
defparam ram40mh_16K_nrnw_inst.INIT_9 = INIT_9;
defparam ram40mh_16K_nrnw_inst.INIT_A = INIT_A;
defparam ram40mh_16K_nrnw_inst.INIT_B = INIT_B;
defparam ram40mh_16K_nrnw_inst.INIT_C = INIT_C;
defparam ram40mh_16K_nrnw_inst.INIT_D = INIT_D;
defparam ram40mh_16K_nrnw_inst.INIT_E = INIT_E;
defparam ram40mh_16K_nrnw_inst.INIT_F = INIT_F;

defparam ram40mh_16K_nrnw_inst.INIT_0 = INIT_0;
defparam ram40mh_16K_nrnw_inst.INIT_1 = INIT_1;
defparam ram40mh_16K_nrnw_inst.INIT_2 = INIT_2;
defparam ram40mh_16K_nrnw_inst.INIT_3 = INIT_3;
defparam ram40mh_16K_nrnw_inst.INIT_4 = INIT_4;
defparam ram40mh_16K_nrnw_inst.INIT_5 = INIT_5;
defparam ram40mh_16K_nrnw_inst.INIT_6 = INIT_6;
defparam ram40mh_16K_nrnw_inst.INIT_7 = INIT_7;
defparam ram40mh_16K_nrnw_inst.INIT_8 = INIT_8;
defparam ram40mh_16K_nrnw_inst.INIT_9 = INIT_9;
defparam ram40mh_16K_nrnw_inst.INIT_A = INIT_A;
defparam ram40mh_16K_nrnw_inst.INIT_B = INIT_B;
defparam ram40mh_16K_nrnw_inst.INIT_C = INIT_C;
defparam ram40mh_16K_nrnw_inst.INIT_D = INIT_D;
defparam ram40mh_16K_nrnw_inst.INIT_E = INIT_E;
defparam ram40mh_16K_nrnw_inst.INIT_F = INIT_F;

`ifdef TIMINGCHECK
specify
   (RCLKN *> RDATA[0]) = (1.0, 1.0);
   (RCLKN *> RDATA[1]) = (1.0, 1.0);
   (RCLKN *> RDATA[2]) = (1.0, 1.0);
   (RCLKN *> RDATA[3]) = (1.0, 1.0);
   (RCLKN *> RDATA[4]) = (1.0, 1.0);
   (RCLKN *> RDATA[5]) = (1.0, 1.0);
   (RCLKN *> RDATA[6]) = (1.0, 1.0);
   (RCLKN *> RDATA[7]) = (1.0, 1.0);
   (RCLKN *> RDATA[8]) = (1.0, 1.0);
   (RCLKN *> RDATA[9]) = (1.0, 1.0);
   (RCLKN *> RDATA[10]) = (1.0, 1.0);
   (RCLKN *> RDATA[11]) = (1.0, 1.0);
   (RCLKN *> RDATA[12]) = (1.0, 1.0);
   (RCLKN *> RDATA[13]) = (1.0, 1.0);
   (RCLKN *> RDATA[14]) = (1.0, 1.0);
   (RCLKN *> RDATA[15]) = (1.0, 1.0);
   $setup(posedge MASK[0], posedge WCLKN, 1.0);
   $setup(negedge MASK[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[0], 1.0);
   $hold(posedge WCLKN, negedge MASK[0], 1.0);
   $setup(posedge MASK[1], posedge WCLKN, 1.0);
   $setup(negedge MASK[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[1], 1.0);
   $hold(posedge WCLKN, negedge MASK[1], 1.0);
   $setup(posedge MASK[2], posedge WCLKN, 1.0);
   $setup(negedge MASK[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[2], 1.0);
   $hold(posedge WCLKN, negedge MASK[2], 1.0);
   $setup(posedge MASK[3], posedge WCLKN, 1.0);
   $setup(negedge MASK[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[3], 1.0);
   $hold(posedge WCLKN, negedge MASK[3], 1.0);
   $setup(posedge MASK[4], posedge WCLKN, 1.0);
   $setup(negedge MASK[4], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[4], 1.0);
   $hold(posedge WCLKN, negedge MASK[4], 1.0);
   $setup(posedge MASK[5], posedge WCLKN, 1.0);
   $setup(negedge MASK[5], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[5], 1.0);
   $hold(posedge WCLKN, negedge MASK[5], 1.0);
   $setup(posedge MASK[6], posedge WCLKN, 1.0);
   $setup(negedge MASK[6], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[6], 1.0);
   $hold(posedge WCLKN, negedge MASK[6], 1.0);
   $setup(posedge MASK[7], posedge WCLKN, 1.0);
   $setup(negedge MASK[7], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[7], 1.0);
   $hold(posedge WCLKN, negedge MASK[7], 1.0);
   $setup(posedge MASK[8], posedge WCLKN, 1.0);
   $setup(negedge MASK[8], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[8], 1.0);
   $hold(posedge WCLKN, negedge MASK[8], 1.0);
   $setup(posedge MASK[9], posedge WCLKN, 1.0);
   $setup(negedge MASK[9], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[9], 1.0);
   $hold(posedge WCLKN, negedge MASK[9], 1.0);
   $setup(posedge MASK[10], posedge WCLKN, 1.0);
   $setup(negedge MASK[10], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[10], 1.0);
   $hold(posedge WCLKN, negedge MASK[10], 1.0);
   $setup(posedge MASK[11], posedge WCLKN, 1.0);
   $setup(negedge MASK[11], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[11], 1.0);
   $hold(posedge WCLKN, negedge MASK[11], 1.0);
   $setup(posedge MASK[12], posedge WCLKN, 1.0);
   $setup(negedge MASK[12], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[12], 1.0);
   $hold(posedge WCLKN, negedge MASK[12], 1.0);
   $setup(posedge MASK[13], posedge WCLKN, 1.0);
   $setup(negedge MASK[13], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[13], 1.0);
   $hold(posedge WCLKN, negedge MASK[13], 1.0);
   $setup(posedge MASK[14], posedge WCLKN, 1.0);
   $setup(negedge MASK[14], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[14], 1.0);
   $hold(posedge WCLKN, negedge MASK[14], 1.0);
   $setup(posedge MASK[15], posedge WCLKN, 1.0);
   $setup(negedge MASK[15], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge MASK[15], 1.0);
   $hold(posedge WCLKN, negedge MASK[15], 1.0);
   $setup(posedge WADDR[0], posedge WCLKN, 1.0);
   $setup(negedge WADDR[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[0], 1.0);
   $hold(posedge WCLKN, negedge WADDR[0], 1.0);
   $setup(posedge WADDR[1], posedge WCLKN, 1.0);
   $setup(negedge WADDR[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[1], 1.0);
   $hold(posedge WCLKN, negedge WADDR[1], 1.0);
   $setup(posedge WADDR[2], posedge WCLKN, 1.0);
   $setup(negedge WADDR[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[2], 1.0);
   $hold(posedge WCLKN, negedge WADDR[2], 1.0);
   $setup(posedge WADDR[3], posedge WCLKN, 1.0);
   $setup(negedge WADDR[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[3], 1.0);
   $hold(posedge WCLKN, negedge WADDR[3], 1.0);
   $setup(posedge WADDR[4], posedge WCLKN, 1.0);
   $setup(negedge WADDR[4], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[4], 1.0);
   $hold(posedge WCLKN, negedge WADDR[4], 1.0);
   $setup(posedge WADDR[5], posedge WCLKN, 1.0);
   $setup(negedge WADDR[5], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[5], 1.0);
   $hold(posedge WCLKN, negedge WADDR[5], 1.0);
   $setup(posedge WADDR[6], posedge WCLKN, 1.0);
   $setup(negedge WADDR[6], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[6], 1.0);
   $hold(posedge WCLKN, negedge WADDR[6], 1.0);
   $setup(posedge WADDR[7], posedge WCLKN, 1.0);
   $setup(negedge WADDR[7], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[7], 1.0);
   $hold(posedge WCLKN, negedge WADDR[7], 1.0);
   $setup(posedge WADDR[8], posedge WCLKN, 1.0);
   $setup(negedge WADDR[8], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[8], 1.0);
   $hold(posedge WCLKN, negedge WADDR[8], 1.0);
   $setup(posedge WADDR[9], posedge WCLKN, 1.0);
   $setup(negedge WADDR[9], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[9], 1.0);
   $hold(posedge WCLKN, negedge WADDR[9], 1.0);
   $setup(posedge WADDR[10], posedge WCLKN, 1.0);
   $setup(negedge WADDR[10], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[10], 1.0);
   $hold(posedge WCLKN, negedge WADDR[10], 1.0);
   $setup(posedge WADDR[11], posedge WCLKN, 1.0);
   $setup(negedge WADDR[11], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[11], 1.0);
   $hold(posedge WCLKN, negedge WADDR[11], 1.0);
   $setup(posedge WADDR[12], posedge WCLKN, 1.0);
   $setup(negedge WADDR[12], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WADDR[12], 1.0);
   $hold(posedge WCLKN, negedge WADDR[12], 1.0);
   $setup(posedge WDATA[0], posedge WCLKN, 1.0);
   $setup(negedge WDATA[0], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[0], 1.0);
   $hold(posedge WCLKN, negedge WDATA[0], 1.0);
   $setup(posedge WDATA[1], posedge WCLKN, 1.0);
   $setup(negedge WDATA[1], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[1], 1.0);
   $hold(posedge WCLKN, negedge WDATA[1], 1.0);
   $setup(posedge WDATA[2], posedge WCLKN, 1.0);
   $setup(negedge WDATA[2], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[2], 1.0);
   $hold(posedge WCLKN, negedge WDATA[2], 1.0);
   $setup(posedge WDATA[3], posedge WCLKN, 1.0);
   $setup(negedge WDATA[3], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[3], 1.0);
   $hold(posedge WCLKN, negedge WDATA[3], 1.0);
   $setup(posedge WDATA[4], posedge WCLKN, 1.0);
   $setup(negedge WDATA[4], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[4], 1.0);
   $hold(posedge WCLKN, negedge WDATA[4], 1.0);
   $setup(posedge WDATA[5], posedge WCLKN, 1.0);
   $setup(negedge WDATA[5], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[5], 1.0);
   $hold(posedge WCLKN, negedge WDATA[5], 1.0);
   $setup(posedge WDATA[6], posedge WCLKN, 1.0);
   $setup(negedge WDATA[6], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[6], 1.0);
   $hold(posedge WCLKN, negedge WDATA[6], 1.0);
   $setup(posedge WDATA[7], posedge WCLKN, 1.0);
   $setup(negedge WDATA[7], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[7], 1.0);
   $hold(posedge WCLKN, negedge WDATA[7], 1.0);
   $setup(posedge WDATA[8], posedge WCLKN, 1.0);
   $setup(negedge WDATA[8], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[8], 1.0);
   $hold(posedge WCLKN, negedge WDATA[8], 1.0);
   $setup(posedge WDATA[9], posedge WCLKN, 1.0);
   $setup(negedge WDATA[9], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[9], 1.0);
   $hold(posedge WCLKN, negedge WDATA[9], 1.0);
   $setup(posedge WDATA[10], posedge WCLKN, 1.0);
   $setup(negedge WDATA[10], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[10], 1.0);
   $hold(posedge WCLKN, negedge WDATA[10], 1.0);
   $setup(posedge WDATA[11], posedge WCLKN, 1.0);
   $setup(negedge WDATA[11], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[11], 1.0);
   $hold(posedge WCLKN, negedge WDATA[11], 1.0);
   $setup(posedge WDATA[12], posedge WCLKN, 1.0);
   $setup(negedge WDATA[12], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[12], 1.0);
   $hold(posedge WCLKN, negedge WDATA[12], 1.0);
   $setup(posedge WDATA[13], posedge WCLKN, 1.0);
   $setup(negedge WDATA[13], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[13], 1.0);
   $hold(posedge WCLKN, negedge WDATA[13], 1.0);
   $setup(posedge WDATA[14], posedge WCLKN, 1.0);
   $setup(negedge WDATA[14], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[14], 1.0);
   $hold(posedge WCLKN, negedge WDATA[14], 1.0);
   $setup(posedge WDATA[15], posedge WCLKN, 1.0);
   $setup(negedge WDATA[15], posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WDATA[15], 1.0);
   $hold(posedge WCLKN, negedge WDATA[15], 1.0);
   $setup(posedge WCLKE, posedge WCLKN, 1.0);
   $setup(negedge WCLKE, posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WCLKE, 1.0);
   $hold(posedge WCLKN, negedge WCLKE, 1.0);
   $setup(posedge WE, posedge WCLKN, 1.0);
   $setup(negedge WE, posedge WCLKN, 1.0);
   $hold(posedge WCLKN, posedge WE, 1.0);
   $hold(posedge WCLKN, negedge WE, 1.0);
   $setup(posedge RADDR[0], posedge RCLKN, 1.0);
   $setup(negedge RADDR[0], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[0], 1.0);
   $hold(posedge RCLKN, negedge RADDR[0], 1.0);
   $setup(posedge RADDR[1], posedge RCLKN, 1.0);
   $setup(negedge RADDR[1], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[1], 1.0);
   $hold(posedge RCLKN, negedge RADDR[1], 1.0);
   $setup(posedge RADDR[2], posedge RCLKN, 1.0);
   $setup(negedge RADDR[2], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[2], 1.0);
   $hold(posedge RCLKN, negedge RADDR[2], 1.0);
   $setup(posedge RADDR[3], posedge RCLKN, 1.0);
   $setup(negedge RADDR[3], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[3], 1.0);
   $hold(posedge RCLKN, negedge RADDR[3], 1.0);
   $setup(posedge RADDR[4], posedge RCLKN, 1.0);
   $setup(negedge RADDR[4], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[4], 1.0);
   $hold(posedge RCLKN, negedge RADDR[4], 1.0);
   $setup(posedge RADDR[5], posedge RCLKN, 1.0);
   $setup(negedge RADDR[5], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[5], 1.0);
   $hold(posedge RCLKN, negedge RADDR[5], 1.0);
   $setup(posedge RADDR[6], posedge RCLKN, 1.0);
   $setup(negedge RADDR[6], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[6], 1.0);
   $hold(posedge RCLKN, negedge RADDR[6], 1.0);
   $setup(posedge RADDR[7], posedge RCLKN, 1.0);
   $setup(negedge RADDR[7], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[7], 1.0);
   $hold(posedge RCLKN, negedge RADDR[7], 1.0);
   $setup(posedge RADDR[8], posedge RCLKN, 1.0);
   $setup(negedge RADDR[8], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[8], 1.0);
   $hold(posedge RCLKN, negedge RADDR[8], 1.0);
   $setup(posedge RADDR[9], posedge RCLKN, 1.0);
   $setup(negedge RADDR[9], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[9], 1.0);
   $hold(posedge RCLKN, negedge RADDR[9], 1.0);
   $setup(posedge RADDR[10], posedge RCLKN, 1.0);
   $setup(negedge RADDR[10], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[10], 1.0);
   $hold(posedge RCLKN, negedge RADDR[10], 1.0);
   $setup(posedge RADDR[11], posedge RCLKN, 1.0);
   $setup(negedge RADDR[11], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[11], 1.0);
   $hold(posedge RCLKN, negedge RADDR[11], 1.0);
   $setup(posedge RADDR[12], posedge RCLKN, 1.0);
   $setup(negedge RADDR[12], posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RADDR[12], 1.0);
   $hold(posedge RCLKN, negedge RADDR[12], 1.0);
   $setup(posedge RCLKE, posedge RCLKN, 1.0);
   $setup(negedge RCLKE, posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RCLKE, 1.0);
   $hold(posedge RCLKN, negedge RCLKE, 1.0);
   $setup(posedge RE, posedge RCLKN, 1.0);
   $setup(negedge RE, posedge RCLKN, 1.0);
   $hold(posedge RCLKN, posedge RE, 1.0);
   $hold(posedge RCLKN, negedge RE, 1.0);
endspecify
`endif

endmodule // SB_RAM40_16KNRNW

// Lightning  IP  // 

//-----------------------------------
// 	---- SB_I2C ----- 
//-----------------------------------

`timescale 1 ns / 1 ps


module SB_I2C (
input  SBCLKI,
input  SBRWI,
input  SBSTBI,
input  SBADRI7,
input  SBADRI6,
input  SBADRI5,
input  SBADRI4,
input  SBADRI3,
input  SBADRI2,
input  SBADRI1,
input  SBADRI0,
input  SBDATI7,
input  SBDATI6,
input  SBDATI5,
input  SBDATI4,
input  SBDATI3,
input  SBDATI2,
input  SBDATI1,
input  SBDATI0,
input  SCLI,
input  SDAI,

output SBDATO7,
output SBDATO6,
output SBDATO5,
output SBDATO4,
output SBDATO3,
output SBDATO2,
output SBDATO1,
output SBDATO0,
output SBACKO,
output I2CIRQ,
output I2CWKUP,
inout SCLO,
output SCLOE,
output SDAO,
output SDAOE);


  parameter I2C_SLAVE_INIT_ADDR = "0b1111100001";
  parameter BUS_ADDR74 = "0b0001";
  // parameter delay50=50000;

wire master, slave;
//reg SDAI_D;

SB_I2C_CORE inst (
 	.SBCLKI(SBCLKI),
 	.SBRWI(SBRWI),
 	.SBSTBI(SBSTBI),
 	.SBADRI7(SBADRI7),
 	.SBADRI6(SBADRI6),
 	.SBADRI5(SBADRI5),
 	.SBADRI4(SBADRI4),
 	.SBADRI3(SBADRI3),
 	.SBADRI2(SBADRI2),
 	.SBADRI1(SBADRI1),
 	.SBADRI0(SBADRI0),
 	.SBDATI7(SBDATI7),
 	.SBDATI6(SBDATI6),
 	.SBDATI5(SBDATI5),
 	.SBDATI4(SBDATI4),
 	.SBDATI3(SBDATI3),
 	.SBDATI2(SBDATI2),
 	.SBDATI1(SBDATI1),
 	.SBDATI0(SBDATI0),
 	.SCLI(SCLI),
 	.SDAI(SDAI),

	.SBDATO7(SBDATO7),
	.SBDATO6(SBDATO6),
	.SBDATO5(SBDATO5),
	.SBDATO4(SBDATO4),
	.SBDATO3(SBDATO3),
	.SBDATO2(SBDATO2),
	.SBDATO1(SBDATO1),
	.SBDATO0(SBDATO0),
	.SBACKO(SBACKO),
	.I2CIRQ(I2CIRQ),
	.I2CWKUP(I2CWKUP),
	.SCLO(SCLO),
	.SCLOE(SCLOE),
	.SDAO(SDAO),
	.SDAOE(SDAOE));
  defparam inst.I2C_SLAVE_INIT_ADDR = I2C_SLAVE_INIT_ADDR;
  defparam inst.BUS_ADDR74 = BUS_ADDR74;

initial begin
	if (BUS_ADDR74!="0b0001" && BUS_ADDR74!="0b0011")
$display ("ID:BUS_ADDR74: should be LLC=0b0001 or LRC=0b0011, otherwise there would be an error ");
end
// always @ (SDAI) 
	// begin
		// SDAI_D <= #delay50 SDAI;
	// end	 
`ifdef TIMINGCHECK

reg NOTIFIER;
specify

   //(SBCLKI *> SCLO) = (1.0, 1.0);

   (SBCLKI *> SBDATO0) = (1.0, 1.0);
   (SBCLKI *> SBDATO1) = (1.0, 1.0);
   (SBCLKI *> SBDATO2) = (1.0, 1.0);
   (SBCLKI *> SBDATO3) = (1.0, 1.0);
   (SBCLKI *> SBDATO4) = (1.0, 1.0);
   (SBCLKI *> SBDATO5) = (1.0, 1.0);
   (SBCLKI *> SBDATO6) = (1.0, 1.0);
   (SBCLKI *> SBDATO7) = (1.0, 1.0);
   (SBCLKI *> SBACKO) = (1.0, 1.0);
   (SBCLKI *> I2CIRQ) = (1.0, 1.0);
   (SBCLKI *> I2CWKUP) = (1.0, 1.0);

    (SCLO *> SDAO) = (1.0, 1.0);
    (SCLO *> SDAOE) = (1.0, 1.0);
    (SCLI *> SDAO) = (1.0, 1.0);
    (SCLI *> SDAOE) = (1.0, 1.0);

   $setup(posedge SBRWI, posedge SBCLKI, 1.0);
   $setup(negedge SBRWI, posedge SBCLKI, 1.0);
   $hold(posedge SBCLKI, posedge SBRWI, 1.0);
   $hold(posedge SBCLKI, negedge SBRWI, 1.0);	 

   $setup(posedge SBSTBI, posedge SBCLKI, 1.0);
   $setup(negedge SBSTBI, posedge SBCLKI, 1.0);
   $hold(posedge SBCLKI, posedge SBSTBI, 1.0);
   $hold(posedge SBCLKI, negedge SBSTBI, 1.0);

   $setup(posedge SBADRI7, posedge SBCLKI, 1.0);
   $setup(negedge SBADRI7, posedge SBCLKI, 1.0);
   $hold(posedge SBCLKI, posedge SBADRI7, 1.0);
   $hold(posedge SBCLKI, negedge SBADRI7, 1.0);

   $setup(posedge SBADRI6, posedge SBCLKI, 1.0);
   $setup(negedge SBADRI6, posedge SBCLKI, 1.0);
   $hold(posedge SBCLKI, posedge SBADRI6, 1.0);
   $hold(posedge SBCLKI, negedge SBADRI6, 1.0);

   $setup(posedge SBADRI5, posedge SBCLKI, 1.0);
   $setup(negedge SBADRI5, posedge SBCLKI, 1.0);
   $hold(posedge SBCLKI, posedge SBADRI5, 1.0);
   $hold(posedge SBCLKI, negedge SBADRI5, 1.0);

   $setup(posedge SBADRI4, posedge SBCLKI, 1.0);
   $setup(negedge SBADRI4, posedge SBCLKI, 1.0);
   $hold(posedge SBCLKI, posedge SBADRI4, 1.0);
   $hold(posedge SBCLKI, negedge SBADRI4, 1.0);

   $setup(posedge SBADRI3, posedge SBCLKI, 1.0);
   $setup(negedge SBADRI3, posedge SBCLKI, 1.0);
   $hold(posedge SBCLKI, posedge SBADRI3, 1.0);
   $hold(posedge SBCLKI, negedge SBADRI3, 1.0);

   $setup(posedge SBADRI2, posedge SBCLKI, 1.0);
   $setup(negedge SBADRI2, posedge SBCLKI, 1.0);
   $hold(posedge SBCLKI, posedge SBADRI2, 1.0);
   $hold(posedge SBCLKI, negedge SBADRI2, 1.0);

   $setup(posedge SBADRI1, posedge SBCLKI, 1.0);
   $setup(negedge SBADRI1, posedge SBCLKI, 1.0);
   $hold(posedge SBCLKI, posedge SBADRI1, 1.0);
   $hold(posedge SBCLKI, negedge SBADRI1, 1.0);

   $setup(posedge SBADRI0, posedge SBCLKI, 1.0);
   $setup(negedge SBADRI0, posedge SBCLKI, 1.0);
   $hold(posedge SBCLKI, posedge SBADRI0, 1.0);
   $hold(posedge SBCLKI, negedge SBADRI0, 1.0);


   $setup(posedge SBDATI7, posedge SBCLKI, 1.0);
   $setup(negedge SBDATI7, posedge SBCLKI, 1.0);
   $hold(posedge SBCLKI, posedge SBDATI7, 1.0);
   $hold(posedge SBCLKI, negedge SBDATI7, 1.0);

   $setup(posedge SBDATI6, posedge SBCLKI, 1.0);
   $setup(negedge SBDATI6, posedge SBCLKI, 1.0);
   $hold(posedge SBCLKI, posedge SBDATI6, 1.0);
   $hold(posedge SBCLKI, negedge SBDATI6, 1.0);

   $setup(posedge SBDATI5, posedge SBCLKI, 1.0);
   $setup(negedge SBDATI5, posedge SBCLKI, 1.0);
   $hold(posedge SBCLKI, posedge SBDATI5, 1.0);
   $hold(posedge SBCLKI, negedge SBDATI5, 1.0);

   $setup(posedge SBDATI4, posedge SBCLKI, 1.0);
   $setup(negedge SBDATI4, posedge SBCLKI, 1.0);
   $hold(posedge SBCLKI, posedge SBDATI4, 1.0);
   $hold(posedge SBCLKI, negedge SBDATI4, 1.0);

   $setup(posedge SBDATI3, posedge SBCLKI, 1.0);
   $setup(negedge SBDATI3, posedge SBCLKI, 1.0);
   $hold(posedge SBCLKI, posedge SBDATI3, 1.0);
   $hold(posedge SBCLKI, negedge SBDATI3, 1.0);

   $setup(posedge SBDATI2, posedge SBCLKI, 1.0);
   $setup(negedge SBDATI2, posedge SBCLKI, 1.0);
   $hold(posedge SBCLKI, posedge SBDATI2, 1.0);
   $hold(posedge SBCLKI, negedge SBDATI2, 1.0);

   $setup(posedge SBDATI1, posedge SBCLKI, 1.0);
   $setup(negedge SBDATI1, posedge SBCLKI, 1.0);
   $hold(posedge SBCLKI, posedge SBDATI1, 1.0);
   $hold(posedge SBCLKI, negedge SBDATI1, 1.0);

   $setup(posedge SBDATI0, posedge SBCLKI, 1.0);
   $setup(negedge SBDATI0, posedge SBCLKI, 1.0);
   $hold(posedge SBCLKI, posedge SBDATI0, 1.0);
   $hold(posedge SBCLKI, negedge SBDATI0, 1.0);

   $setuphold(posedge SCLO, posedge SDAI, 1.0, 1.0, NOTIFIER);
   $setuphold(posedge SCLO, negedge SDAI, 1.0, 1.0, NOTIFIER);

   $setuphold(posedge SCLI, posedge SDAI, 1.0, 1.0, NOTIFIER);
   $setuphold(posedge SCLI, negedge SDAI, 1.0, 1.0, NOTIFIER);

endspecify
`endif


endmodule



//------------------------------------------
//     ---- SB_SPI  ---- 
//------------------------------------------

`timescale 1 ns / 1 ps

module SB_SPI (
input  SBCLKI,
input  SBRWI,				   
input  SBSTBI,
input  SBADRI7,
input  SBADRI6,
input  SBADRI5,
input  SBADRI4,
input  SBADRI3,
input  SBADRI2,
input  SBADRI1,
input  SBADRI0,
input  SBDATI7,
input  SBDATI6,
input  SBDATI5,
input  SBDATI4,
input  SBDATI3,
input  SBDATI2,
input  SBDATI1,
input  SBDATI0,
input  MI,
input  SI,
input  SCKI,
input  SCSNI,

output SBDATO7,
output SBDATO6,
output SBDATO5,
output SBDATO4,
output SBDATO3,
output SBDATO2,
output SBDATO1,
output SBDATO0,
output SBACKO,
output SPIIRQ,
output SPIWKUP,
output SO,
output SOE,
output MO,
output MOE,
inout SCKO,
output SCKOE,
output MCSNO3,
output MCSNO2,
output MCSNO1,
output MCSNO0,
output MCSNOE3,
output MCSNOE2,
output MCSNOE1,
output MCSNOE0);

parameter BUS_ADDR74 = "0b0000";

SB_SPI_CORE inst (
	.SBCLKI(SBCLKI),
	.SBRWI(SBRWI),
	.SBSTBI(SBSTBI),
	.SBADRI7(SBADRI7),
	.SBADRI6(SBADRI6),
	.SBADRI5(SBADRI5),
	.SBADRI4(SBADRI4),
	.SBADRI3(SBADRI3),
	.SBADRI2(SBADRI2),
	.SBADRI1(SBADRI1),
	.SBADRI0(SBADRI0),
	.SBDATI7(SBDATI7),
	.SBDATI6(SBDATI6),
	.SBDATI5(SBDATI5),
	.SBDATI4(SBDATI4),
	.SBDATI3(SBDATI3),
	.SBDATI2(SBDATI2),
	.SBDATI1(SBDATI1),
	.SBDATI0(SBDATI0),
	.MI(MI),
	.SI(SI),
	.SCKI(SCKI),
	.SCSNI(SCSNI),

	.SBDATO7(SBDATO7),
	.SBDATO6(SBDATO6),
	.SBDATO5(SBDATO5),
	.SBDATO4(SBDATO4),
	.SBDATO3(SBDATO3),
	.SBDATO2(SBDATO2),
	.SBDATO1(SBDATO1),
	.SBDATO0(SBDATO0),
	.SBACKO(SBACKO),
	.SPIIRQ(SPIIRQ),
	.SPIWKUP(SPIWKUP),
	.SO(SO),
	.SOE(SOE),
	.MO(MO),
	.MOE(MOE),
	.SCKO(SCKO),
	.SCKOE(SCKOE),
	.MCSNO3(MCSNO3),
	.MCSNO2(MCSNO2),
	.MCSNO1(MCSNO1),
	.MCSNO0(MCSNO0),
	.MCSNOE3(MCSNOE3),
	.MCSNOE2(MCSNOE2),
	.MCSNOE1(MCSNOE1),
	.MCSNOE0(MCSNOE0));
defparam inst.BUS_ADDR74 = BUS_ADDR74;

initial begin
	if (BUS_ADDR74!="0b0000" && BUS_ADDR74!="0b0010")
$display ("ID:BUS_ADDR74: should be LLC=0b0000 or LRC=0b0010, otherwise there would be an error ");
end

`ifdef TIMINGCHECK

reg NOTIFIER;

specify

	//(SBCLKI *> SCKO) = (1.0, 1.0);

	(SBCLKI *> SBDATO0) = (1.0, 1.0);
	(SBCLKI *> SBDATO1) = (1.0, 1.0);
	(SBCLKI *> SBDATO2) = (1.0, 1.0);
	(SBCLKI *> SBDATO3) = (1.0, 1.0);
	(SBCLKI *> SBDATO4) = (1.0, 1.0);
	(SBCLKI *> SBDATO5) = (1.0, 1.0);
	(SBCLKI *> SBDATO6) = (1.0, 1.0);
	(SBCLKI *> SBDATO7) = (1.0, 1.0);
	(SBCLKI *> SBACKO) = (1.0, 1.0);
	(SBCLKI *> SPIIRQ) = (1.0, 1.0);
	(SBCLKI *> SPIWKUP) = (1.0, 1.0);

	(SCKO *> MO) = (1.0, 1.0);
	(SCKO *> MOE) = (1.0, 1.0);
	(SCKO *> MCSNO3) = (1.0, 1.0);
	(SCKO *> MCSNO2) = (1.0, 1.0);
	(SCKO *> MCSNO1) = (1.0, 1.0);
	(SCKO *> MCSNO0) = (1.0, 1.0);
	(SCKO *> MCSNOE3) = (1.0, 1.0);
	(SCKO *> MCSNOE2) = (1.0, 1.0);
	(SCKO *> MCSNOE1) = (1.0, 1.0);
	(SCKO *> MCSNOE0) = (1.0, 1.0);

       	(SCKI *> SO) = (1.0, 1.0);
       	(SCKI *> SOE) = (1.0, 1.0);	  
		   
	
//	$setup(posedge 	SBRWI, negedge SBCLKI, 1.0);
//	$setup(negedge 	SBRWI, negedge SBCLKI, 1.0); 
	$setup(posedge 	SBRWI, posedge SBCLKI, 1.0);
	$setup(negedge 	SBRWI, posedge SBCLKI, 1.0); 
	$hold(posedge SBCLKI, posedge SBRWI, 1.0);
	$hold(posedge SBCLKI, negedge SBRWI, 1.0);

	$setup(posedge 	SBSTBI, posedge SBCLKI, 1.0);
	$setup(negedge 	SBSTBI, posedge SBCLKI, 1.0);
	$hold(posedge SBCLKI, posedge SBSTBI, 1.0);
	$hold(posedge SBCLKI, negedge SBSTBI, 1.0);
	   
	$setup(posedge 	SBADRI7, posedge SBCLKI, 1.0);
	$setup(negedge 	SBADRI7, posedge SBCLKI, 1.0);
	$hold(posedge SBCLKI, posedge SBADRI7, 1.0);
	$hold(posedge SBCLKI, negedge SBADRI7, 1.0);
	$setup(posedge 	SBADRI6, posedge SBCLKI, 1.0);
	$setup(negedge 	SBADRI6, posedge SBCLKI, 1.0);
	$hold(posedge SBCLKI, posedge SBADRI6, 1.0);
	$hold(posedge SBCLKI, negedge SBADRI6, 1.0);
	$setup(posedge 	SBADRI5, posedge SBCLKI, 1.0);
	$setup(negedge 	SBADRI5, posedge SBCLKI, 1.0);
	$hold(posedge SBCLKI, posedge SBADRI5, 1.0);
	$hold(posedge SBCLKI, negedge SBADRI5, 1.0);
	$setup(posedge 	SBADRI4, posedge SBCLKI, 1.0);
	$setup(negedge 	SBADRI4, posedge SBCLKI, 1.0);
	$hold(posedge SBCLKI, posedge SBADRI4, 1.0);
	$hold(posedge SBCLKI, negedge SBADRI4, 1.0);
	$setup(posedge 	SBADRI3, posedge SBCLKI, 1.0);
	$setup(negedge 	SBADRI3, posedge SBCLKI, 1.0);
	$hold(posedge SBCLKI, posedge SBADRI3, 1.0);
	$hold(posedge SBCLKI, negedge SBADRI3, 1.0);
	$setup(posedge 	SBADRI2, posedge SBCLKI, 1.0);
	$setup(negedge 	SBADRI2, posedge SBCLKI, 1.0);
	$hold(posedge SBCLKI, posedge SBADRI2, 1.0);
	$hold(posedge SBCLKI, negedge SBADRI2, 1.0);
	$setup(posedge 	SBADRI1, posedge SBCLKI, 1.0);
	$setup(negedge 	SBADRI1, posedge SBCLKI, 1.0);
	$hold(posedge SBCLKI, posedge SBADRI1, 1.0);
	$hold(posedge SBCLKI, negedge SBADRI1, 1.0);
	$setup(posedge 	SBADRI0, posedge SBCLKI, 1.0);
	$setup(negedge 	SBADRI0, posedge SBCLKI, 1.0);
	$hold(posedge SBCLKI, posedge SBADRI0, 1.0);
	$hold(posedge SBCLKI, negedge SBADRI0, 1.0);

	$setup(posedge 	SBDATI7, posedge SBCLKI, 1.0);
	$setup(negedge 	SBDATI7, posedge SBCLKI, 1.0);
	$hold(posedge SBCLKI, posedge SBDATI7, 1.0);
	$hold(posedge SBCLKI, negedge SBDATI7, 1.0);
	$setup(posedge 	SBDATI6, posedge SBCLKI, 1.0);
	$setup(negedge 	SBDATI6, posedge SBCLKI, 1.0);
	$hold(posedge SBCLKI, posedge SBDATI6, 1.0);
	$hold(posedge SBCLKI, negedge SBDATI6, 1.0);
	$setup(posedge 	SBDATI5, posedge SBCLKI, 1.0);
	$setup(negedge 	SBDATI5, posedge SBCLKI, 1.0);
	$hold(posedge SBCLKI, posedge SBDATI5, 1.0);
	$hold(posedge SBCLKI, negedge SBDATI5, 1.0);
	$setup(posedge 	SBDATI4, posedge SBCLKI, 1.0);
	$setup(negedge 	SBDATI4, posedge SBCLKI, 1.0);
	$hold(posedge SBCLKI, posedge SBDATI4, 1.0);
	$hold(posedge SBCLKI, negedge SBDATI4, 1.0);
	$setup(posedge 	SBDATI3, posedge SBCLKI, 1.0);
	$setup(negedge 	SBDATI3, posedge SBCLKI, 1.0);
	$hold(posedge SBCLKI, posedge SBDATI3, 1.0);
	$hold(posedge SBCLKI, negedge SBDATI3, 1.0);
	$setup(posedge 	SBDATI2, posedge SBCLKI, 1.0);
	$setup(negedge 	SBDATI2, posedge SBCLKI, 1.0);
	$hold(posedge SBCLKI, posedge SBDATI2, 1.0);
	$hold(posedge SBCLKI, negedge SBDATI2, 1.0);
	$setup(posedge 	SBDATI1, posedge SBCLKI, 1.0);
	$setup(negedge 	SBDATI1, posedge SBCLKI, 1.0);
	$hold(posedge SBCLKI, posedge SBDATI1, 1.0);
	$hold(posedge SBCLKI, negedge SBDATI1, 1.0);
	$setup(posedge 	SBDATI0, posedge SBCLKI, 1.0);
	$setup(negedge 	SBDATI0, posedge SBCLKI, 1.0);
	$hold(posedge SBCLKI, posedge SBDATI0, 1.0);
	$hold(posedge SBCLKI, negedge SBDATI0, 1.0);

	$setuphold(posedge SCKO, posedge 	MI, 1.0, 1.0, NOTIFIER);
	$setuphold(posedge SCKO, negedge 	MI, 1.0, 1.0, NOTIFIER);

	$setuphold(posedge SCKI, posedge SI, 1.0, 1.0, NOTIFIER);
	$setuphold(posedge SCKI, negedge SI, 1.0, 1.0, NOTIFIER);

	$setuphold(posedge SCKI, posedge SCSNI, 1.0, 1.0, NOTIFIER);
	$setuphold(posedge SCKI, negedge SCSNI, 1.0, 1.0, NOTIFIER);  
		/////////////////////added/////////////////	
	 
	$setuphold(negedge SCKO, posedge 	MI, 1.0, 1.0, NOTIFIER);
	$setuphold(negedge SCKO, negedge 	MI, 1.0, 1.0, NOTIFIER);

	$setuphold(negedge SCKI, posedge SI, 1.0, 1.0, NOTIFIER);
	$setuphold(negedge SCKI, negedge SI, 1.0, 1.0, NOTIFIER);

	$setuphold(negedge SCKI, posedge SCSNI, 1.0, 1.0, NOTIFIER);
	$setuphold(negedge SCKI, negedge SCSNI, 1.0, 1.0, NOTIFIER); 

endspecify	  
`endif
endmodule
//--------------------------------------
//    ---  SB_HSOSC ----- 
//-------------------------------------- 

`timescale 1 ns / 1 ps
module SB_HSOSC (input ENACLKM, output CLKM);  

SB_HSOSC_CORE inst(
	.ENACLKM(ENACLKM),
	.CLKM(CLKM));

`ifdef TIMINGCHECK
specify

   (ENACLKM *> CLKM) = (1.0, 1.0);

endspecify
`endif

endmodule

//--------------------------------------
// ----  SB_LSOSC ------ 
//--------------------------------------

`timescale 1 ns / 1 ps

module SB_LSOSC (input ENACLKK, output CLKK);

SB_LSOSC_CORE inst(
	.ENACLKK(ENACLKK),
	.CLKK(CLKK));  

`ifdef TIMINGCHECK
specify

   (ENACLKK *> CLKK) = (1.0, 1.0);

endspecify
`endif

endmodule

//--------------------------------------
// ----  SB_LFOSC ------ 
//--------------------------------------


`timescale 1ps/1ps
module 	 SB_LFOSC ( CLKLFEN, CLKLFPU,  CLKLF);	 
input CLKLFEN, CLKLFPU;
output CLKLF;	
SB_LFOSC_CORE OSCInst1 ( 
.CLKLF_EN(CLKLFEN), 
.CLKLF_PU(CLKLFPU),
.CLKLF(CLKLF) 
) /* synthesis ROUTE_THROUGH_FABRIC= 0 */;

`ifdef TIMINGCHECK
specify

	//(CLKLFEN *> CLKLF) = (1.0, 1.0);
	(CLKLFPU *> CLKLF) = (1.0, 1.0);
endspecify
`endif

endmodule 

//--------------------------------------
// ----  SB_HFOSC ------ 
//--------------------------------------
`timescale 1ps/1ps
module SB_HFOSC  ( CLKHFPU,CLKHFEN, CLKHF);	
	input CLKHFPU,CLKHFEN;
	output  CLKHF;	
	parameter CLKHF_DIV = "0b00";
SB_HFOSC_CORE OSCInst0( 
.CLKHF_EN(CLKHFEN), 
.CLKHF_PU(CLKHFPU),
.CLKHF(CLKHF) 
) /* synthesis ROUTE_THROUGH_FABRIC= 0 */;
defparam OSCInst0.CLKHF_DIV = CLKHF_DIV;

`ifdef TIMINGCHECK
specify

   (CLKHFPU *> CLKHF) = (1.0, 1.0);
 //  (CLKHFEN *> CLKHF) = (1.0, 1.0);

endspecify
`endif

endmodule 

//--------------------------------------
// ----  SB_IR_DRV ------ 
//--------------------------------------
`timescale 1ps/1ps
module SB_IR_DRV (IRLEDEN,IRPWM,IRPU,IRLED);

input IRLEDEN,IRPWM,IRPU ;
output IRLED;	  

parameter IR_CURRENT = "0b0000000000"; 
SB_IR_DRV_CORE inst (.IRLED_EN(IRLEDEN),.IR_PWM(IRPWM),.IR_PU(IRPU),.IRLED(IRLED));
defparam inst.IR_CURRENT=IR_CURRENT;

`ifdef TIMINGCHECK
specify

   (IRPWM *> IRLED) = (1.0, 1.0);

endspecify
`endif

endmodule
//--------------------------------------
// ----  SB_RGB_DRV ------ 
//--------------------------------------
`timescale 1ps/1ps
module SB_RGB_DRV (RGBLEDEN,RGB0PWM, RGB1PWM ,RGB2PWM, RGBPU, RGB0, RGB1, RGB2 );
input  RGBLEDEN,RGB0PWM, RGB1PWM ,RGB2PWM, RGBPU;
output   RGB0, RGB1, RGB2; 
parameter RGB0_CURRENT = "0b000000";
parameter RGB1_CURRENT = "0b000000";
parameter RGB2_CURRENT = "0b000000";
SB_RGB_DRV_CORE inst (.RGBLED_EN(RGBLEDEN ),.RGB0_PWM( RGB0PWM), .RGB1_PWM (RGB1PWM ),.RGB2_PWM(RGB2PWM ), .RGB_PU( RGBPU), .RGB0( RGB0), .RGB1( RGB1), .RGB2(RGB2));
defparam inst.RGB0_CURRENT= RGB0_CURRENT;
defparam inst.RGB1_CURRENT= RGB1_CURRENT;
defparam inst.RGB2_CURRENT= RGB2_CURRENT;	

`ifdef TIMINGCHECK
specify

   (RGB0PWM *> RGB0) = (1.0, 1.0);
   (RGB1PWM *> RGB1) = (1.0, 1.0);
   (RGB2PWM *> RGB2) = (1.0, 1.0);

endspecify
`endif

endmodule

//--------------------------------------
// ----  LED_DRV_CUR ------ 
//--------------------------------------
`timescale 1ps/1ps
module SB_LED_DRV_CUR  ( EN, LEDPU);
input EN;
output LEDPU;

wire powerup;

   assign powerup = (EN === 1'b1) ? 1'b0 : 1'b1; //Constant current source
   buf (LEDPU, powerup) ;

`ifdef TIMINGCHECK
specify

   (EN *> LEDPU) = (1.0, 1.0);

endspecify
`endif
endmodule
//-------------------------------------
// ----  SB_LEDD_IP ------ 
//--------------------------------------
`timescale 1ps/1ps
module SB_LEDD_IP ( LEDDCS,LEDDCLK,LEDDDAT7,LEDDDAT6,LEDDDAT5,LEDDDAT4,
	LEDDDAT3,LEDDDAT2,LEDDDAT1,LEDDDAT0,LEDDADDR3,LEDDADDR2,LEDDADDR1,
	LEDDADDR0,LEDDDEN,LEDDEXE,LEDDRST,PWMOUT0,PWMOUT1,PWMOUT2,LEDDON);	 
	
	input 	LEDDCS,LEDDCLK,LEDDDAT7,LEDDDAT6,LEDDDAT5,LEDDDAT4,LEDDDAT3,LEDDDAT2,
			LEDDDAT1,LEDDDAT0,LEDDADDR3,LEDDADDR2,LEDDADDR1,LEDDADDR0,LEDDDEN,LEDDEXE,LEDDRST; 
	output  PWMOUT0,PWMOUT1,PWMOUT2,LEDDON;
	
	wire LEDDCS, LEDDCLK,LEDDDAT7,LEDDDAT6,LEDDDAT5,LEDDDAT4,LEDDDAT3,LEDDDAT2, LEDDDAT1,LEDDDAT0,LEDDADDR3,LEDDADDR2,LEDDADDR1,LEDDADDR0,LEDDDEN,LEDDEXE,LEDDRST; 
	wire PWMOUT0,PWMOUT1,PWMOUT2,LEDDON;
	wire [7:0]  sb_ledd_dat={LEDDDAT7,LEDDDAT6,LEDDDAT5, LEDDDAT4,LEDDDAT3,LEDDDAT2,LEDDDAT1,LEDDDAT0};
	wire [3:0]	sb_ledd_adr={LEDDADDR3,LEDDADDR2,LEDDADDR1,LEDDADDR0};
	reg NOTIFIER;
	reg ledd_rst_async;
	initial
begin
   ledd_rst_async = 1'b1;
#100
   ledd_rst_async = 1'b0;
end
	ledd_ip  ledd_ip_inst
	(
	.pwm_out_r(PWMOUT0),
	.pwm_out_g(PWMOUT1), 
	.pwm_out_b(PWMOUT2), 
	.ledd_on(LEDDON),
	.ledd_rst_async(ledd_rst_async), 
	.ledd_clk(LEDDCLK), 
	.ledd_cs(LEDDCS), 
	.ledd_den(LEDDDEN), 
	.ledd_adr(sb_ledd_adr), 
	.ledd_dat(sb_ledd_dat),
    .ledd_exe(LEDDEXE)
   );
   
   `ifdef TIMINGCHECK
specify


	(LEDDCLK*>PWMOUT0) = (1.0, 1.0);
	(LEDDCLK*>PWMOUT1) = (1.0, 1.0);
	(LEDDCLK*>PWMOUT2) = (1.0, 1.0);
	(LEDDCLK*>LEDDON) = (1.0, 1.0);	 
   	$setup(posedge LEDDCS, posedge LEDDCLK,  1.0);  
	$setup(negedge LEDDCS, posedge LEDDCLK,  1.0); 
	$hold(posedge LEDDCLK, posedge LEDDCS,  1.0);
	$hold(posedge LEDDCLK, negedge LEDDCS,  1.0); 
	$setup(posedge LEDDDEN, posedge LEDDCLK,  1.0);  
	$setup(negedge LEDDDEN, posedge LEDDCLK,  1.0); 
	$hold(posedge LEDDCLK, posedge LEDDDEN,  1.0);
	$hold(posedge LEDDCLK, negedge LEDDDEN,  1.0);
	$setup(posedge LEDDEXE, posedge LEDDCLK,  1.0);  
	$setup(negedge LEDDEXE, posedge LEDDCLK,  1.0); 
	$hold(posedge LEDDCLK, posedge LEDDEXE,  1.0);
	$hold(posedge LEDDCLK, negedge LEDDEXE,  1.0);
	$setup(posedge LEDDADDR0, posedge LEDDCLK,  1.0);  
	$setup(negedge LEDDADDR0, posedge LEDDCLK,  1.0); 
	$hold(posedge LEDDCLK, posedge LEDDADDR0,  1.0);
	$hold(posedge LEDDCLK, negedge LEDDADDR0,  1.0);
	$setup(posedge LEDDADDR1, posedge LEDDCLK,  1.0);  
	$setup(negedge LEDDADDR1, posedge LEDDCLK,  1.0); 
	$hold(posedge LEDDCLK, posedge LEDDADDR1,  1.0);
	$hold(posedge LEDDCLK, negedge LEDDADDR1,  1.0);
	$setup(posedge LEDDADDR2, posedge LEDDCLK,  1.0);  
	$setup(negedge LEDDADDR2, posedge LEDDCLK,  1.0); 
	$hold(posedge LEDDCLK, posedge LEDDADDR2,  1.0);
	$hold(posedge LEDDCLK, negedge LEDDADDR2,  1.0);
	$setup(posedge LEDDADDR3, posedge LEDDCLK,  1.0);  
	$setup(negedge LEDDADDR3, posedge LEDDCLK,  1.0); 
	$hold(posedge LEDDCLK, posedge LEDDADDR3,  1.0);
	$hold(posedge LEDDCLK, negedge LEDDADDR3,  1.0);

	$setup(posedge LEDDDAT0, posedge LEDDCLK,  1.0);  
	$setup(negedge LEDDDAT0, posedge LEDDCLK,  1.0); 
	$hold(posedge LEDDCLK, posedge LEDDDAT0,  1.0);
	$hold(posedge LEDDCLK, negedge LEDDDAT0,  1.0);
	$setup(posedge LEDDDAT1, posedge LEDDCLK,  1.0);  
	$setup(negedge LEDDDAT1, posedge LEDDCLK,  1.0); 
	$hold(posedge LEDDCLK, posedge LEDDDAT1,  1.0);
	$hold(posedge LEDDCLK, negedge LEDDDAT1,  1.0);
	$setup(posedge LEDDDAT2, posedge LEDDCLK,  1.0);  
	$setup(negedge LEDDDAT2, posedge LEDDCLK,  1.0); 
	$hold(posedge LEDDCLK, posedge LEDDDAT2,  1.0);
	$hold(posedge LEDDCLK, negedge LEDDDAT2,  1.0);
	$setup(posedge LEDDDAT3, posedge LEDDCLK,  1.0);  
	$setup(negedge LEDDDAT3, posedge LEDDCLK,  1.0); 
	$hold(posedge LEDDCLK, posedge LEDDDAT3,  1.0);
	$hold(posedge LEDDCLK, negedge LEDDDAT3,  1.0);
	$setup(posedge LEDDDAT4, posedge LEDDCLK,  1.0);  
	$setup(negedge LEDDDAT4, posedge LEDDCLK,  1.0); 
	$hold(posedge LEDDCLK, posedge LEDDDAT4,  1.0);
	$hold(posedge LEDDCLK, negedge LEDDDAT4,  1.0);
	$setup(posedge LEDDDAT5, posedge LEDDCLK,  1.0);  
	$setup(negedge LEDDDAT5, posedge LEDDCLK,  1.0); 
	$hold(posedge LEDDCLK, posedge LEDDDAT5,  1.0);
	$hold(posedge LEDDCLK, negedge LEDDDAT5,  1.0);
	$setup(posedge LEDDDAT6, posedge LEDDCLK,  1.0);  
	$setup(negedge LEDDDAT6, posedge LEDDCLK,  1.0); 
	$hold(posedge LEDDCLK, posedge LEDDDAT6,  1.0);
	$hold(posedge LEDDCLK, negedge LEDDDAT6,  1.0);
	$setup(posedge LEDDDAT7, posedge LEDDCLK,  1.0);  
	$setup(negedge LEDDDAT7, posedge LEDDCLK,  1.0); 
	$hold(posedge LEDDCLK, posedge LEDDDAT7,  1.0);
	$hold(posedge LEDDCLK, negedge LEDDDAT7,  1.0);

		 endspecify
`endif

   
endmodule


//--------------------------------------
// ----  SB_IO_OD ------ 
//--------------------------------------
`timescale 1ps/1ps

module SB_IO_OD (
	PACKAGEPIN, 
	LATCHINPUTVALUE, 
	CLOCKENABLE, 
	INPUTCLK, 
	OUTPUTCLK, 
	OUTPUTENABLE, 
	DOUT1, 
	DOUT0, 
	DIN1, 
	DIN0
 );

parameter PIN_TYPE			= 6'b000000;	  // The default is set to report IO macros that do not define what IO type is used. 
//parameter PULLUP = 1'b0; // by default the IO will have NO pullup, this parameter is used only on bank 0, 1, and 2. Will be ignored when it is placed at bank 3
parameter NEG_TRIGGER = 1'b0; // specify the polarity of all FFs in the IO to be falling edge when NEG_TRIGGER = 1, default is rising edge
//parameter IO_STANDARD = "SB_LVCMOS"; // more standards are supported in bank 3 only: SB_SSTL2_CLASS_2, SB_SSTL2_CLASS_1, SB_SSTL18_FULL, SB_SSTL18_HALF
						 // SB_MDDR10, SB_MDDR8, SB_MDDR4, SB_MDDR2

input DOUT1;  		// Input output 1
input DOUT0;  		// Input output 0

input CLOCKENABLE;    		// Clock enables NEW - common to in/out clocks

output DIN1;    		// Output input 1
output DIN0;    		// Output input 0

input OUTPUTENABLE;   		// Ouput-Enable 
input LATCHINPUTVALUE;    		// Input control
input INPUTCLK;   		// Input clock
input OUTPUTCLK;  		// Output clock

inout 	PACKAGEPIN; 		//' User's package pin - 'PAD' output

//------------- Main Body of verilog ----------------------------------------------------
wire inclk_, outclk_;
wire inclk, outclk;
reg INCLKE_sync, OUTCLKE_sync; 

assign (weak0, weak1) CLOCKENABLE =1'b1 ;
assign (weak0, weak1) DOUT0	  =1'b0 ;
assign (weak0, weak1) DOUT1 	  =1'b0 ;
assign inclk_ = (INPUTCLK ^ NEG_TRIGGER); // change the input clock phase
assign outclk_ = (OUTPUTCLK ^ NEG_TRIGGER); // change the output clock phase
//assign inclk = (inclk_ & CLOCK_ENABLE);
//assign outclk = (outclk_ & CLOCK_ENABLE);

//////// CLKEN sync ///////
always@(inclk_ or CLOCKENABLE)
begin 
    if(~inclk_)
	INCLKE_sync = CLOCKENABLE; 
end

always@(outclk_ or CLOCKENABLE)
begin 
   if(~outclk_) 	
	OUTCLKE_sync = CLOCKENABLE; 
end

assign inclk = (inclk_ & INCLKE_sync);
assign outclk = (outclk_ & OUTCLKE_sync);

wire bs_en;   //Boundary scan enable
wire shift;   //Boundary scan shift
wire tclk;    //Boundary scan clock
wire update;  //Boundary scan update
wire sdi;     //Boundary scan serial data in
wire mode;    //Boundary scan mode
wire hiz_b;   //Boundary scan tristate control
wire sdo;     //Boundary scan serial data out

//wire rstio; disabled as this a power on only signal   	//Normal Input reset
assign  bs_en = 1'b0;	//Boundary scan enable
assign  shift = 1'b0;	//Boundary scan shift
assign  tclk = 1'b0;	//Boundary scan clock
assign  update = 1'b0;	//Boundary scan update
assign  sdi = 1'b0;	//Boundary scan serial data in
assign  mode = 1'b0;	//Boundary scan mode
assign  hiz_b = 1'b1;	//Boundary scan Tristate control
  
wire padoen, padout, padin;
assign PACKAGEPIN = ((~padoen) && (~padout)) ? 1'b0 : 1'bz;
assign padin = PACKAGEPIN ;


//parameter Pin_Type  MUST be defined when instantiated
wire hold, oepin;							  // The required package pin type must be set when io_macro is instantiated.
assign hold = LATCHINPUTVALUE;
assign oepin = OUTPUTENABLE;
 
 preio_physical preiophysical_i (	//original names unchanged
 	.hold(hold),
	.rstio(1'b0),			//Disabled as this is power on only.
	.bs_en(bs_en),
	.shift(shift),
	.tclk(tclk),
	.inclk(inclk),
	.outclk(outclk),
	.update(update),
	.oepin(oepin),
	.sdi(sdi),
	.mode(mode),
	.hiz_b(hiz_b),
	.sdo(sdo),
	.dout1(DIN1),
	.dout0(DIN0),
	.ddr1(DOUT1),
	.ddr0(DOUT0),
	.padin(padin),
	.padout(padout),
	.padoen(padoen),
	.cbit(PIN_TYPE)
	);
	`ifdef TIMINGCHECK
specify
   (PACKAGEPIN *> DIN0) = (1.0, 1.0);
   (PACKAGEPIN *> DIN1) = (1.0, 1.0);
   (INPUTCLK *> DIN0) = (1.0, 1.0);
   (INPUTCLK *> DIN1) = (1.0, 1.0);
   (DOUT0 *> PACKAGEPIN) = (1.0, 1.0);
   (DOUT1 *> PACKAGEPIN) = (1.0, 1.0);
   (OUTPUTENABLE *> PACKAGEPIN) = (1.0, 1.0);
   (INPUTCLK *> PACKAGEPIN) = (1.0, 1.0);
   (OUTPUTCLK *> PACKAGEPIN) = (1.0, 1.0);
   (LATCHINPUTVALUE *> DIN0) = (1.0, 1.0);
   (LATCHINPUTVALUE *> DIN1) = (1.0, 1.0);
   $setup(posedge CLOCKENABLE, posedge INPUTCLK, 1.0);
   $setup(negedge CLOCKENABLE, posedge INPUTCLK, 1.0);
   $hold(posedge INPUTCLK, posedge CLOCKENABLE, 1.0);
   $hold(posedge INPUTCLK, negedge CLOCKENABLE, 1.0);
   $setup(posedge PACKAGEPIN, posedge INPUTCLK, 1.0);
   $setup(negedge PACKAGEPIN, posedge INPUTCLK, 1.0);
   $hold(posedge INPUTCLK, posedge PACKAGEPIN, 1.0);
   $hold(posedge INPUTCLK, negedge PACKAGEPIN, 1.0);
   $setup(posedge PACKAGEPIN, negedge INPUTCLK, 1.0);
   $setup(negedge PACKAGEPIN, negedge INPUTCLK, 1.0);
   $hold(negedge INPUTCLK, posedge PACKAGEPIN, 1.0);
   $hold(negedge INPUTCLK, negedge PACKAGEPIN, 1.0);
   $setup(posedge CLOCKENABLE, posedge OUTPUTCLK, 1.0);
   $setup(negedge CLOCKENABLE, posedge OUTPUTCLK, 1.0);
   $hold(posedge OUTPUTCLK, posedge CLOCKENABLE, 1.0);
   $hold(posedge OUTPUTCLK, negedge CLOCKENABLE, 1.0);
   $setup(posedge PACKAGEPIN, posedge OUTPUTCLK, 1.0);
   $setup(negedge PACKAGEPIN, posedge OUTPUTCLK, 1.0);
   $hold(posedge OUTPUTCLK, posedge PACKAGEPIN, 1.0);
   $hold(posedge OUTPUTCLK, negedge PACKAGEPIN, 1.0);
   $setup(posedge DOUT0, posedge OUTPUTCLK, 1.0);
   $setup(negedge DOUT0, posedge OUTPUTCLK, 1.0);
   $hold(posedge OUTPUTCLK, posedge DOUT0, 1.0);
   $hold(posedge OUTPUTCLK, negedge DOUT0, 1.0);
   $setup(posedge DOUT1, posedge OUTPUTCLK, 1.0);
   $setup(negedge DOUT1, posedge OUTPUTCLK, 1.0);
   $hold(posedge OUTPUTCLK, posedge DOUT1, 1.0);
   $hold(posedge OUTPUTCLK, negedge DOUT1, 1.0);
   $setup(posedge DOUT1, negedge OUTPUTCLK, 1.0);
   $setup(negedge DOUT1, negedge OUTPUTCLK, 1.0);
   $hold(negedge OUTPUTCLK, posedge DOUT1, 1.0);
   $hold(negedge OUTPUTCLK, negedge DOUT1, 1.0);
   $setup(posedge DOUT0, posedge OUTPUTCLK, 1.0);
   $setup(negedge DOUT0, posedge OUTPUTCLK, 1.0);
   $hold(posedge OUTPUTCLK, posedge DOUT0, 1.0);
   $hold(posedge OUTPUTCLK, negedge DOUT0, 1.0);
   $setup(posedge OUTPUTENABLE, posedge OUTPUTCLK, 1.0);
   $setup(negedge OUTPUTENABLE, posedge OUTPUTCLK, 1.0);
   $hold(posedge OUTPUTCLK, posedge OUTPUTENABLE, 1.0);
   $hold(posedge OUTPUTCLK, negedge OUTPUTENABLE, 1.0);

endspecify
`endif
endmodule

//--------------------------------------
// ----  SB_RGBA_DRV ------ 
//--------------------------------------
`timescale 1ps/1ps

module SB_RGBA_DRV(RGB0, RGB0PWM, RGB1, RGB1PWM, RGB2, RGB2PWM, CURREN, RGBLEDEN); 

// *** Input to UUT ***
input            RGB0PWM;
 input            RGB1PWM;
 input            RGB2PWM;
 input            CURREN;
 input            RGBLEDEN;

// *** Inouts to UUT ***

// *** Outputs from UUT ***
output            RGB0;
 output            RGB1;
 output            RGB2;

parameter          CURRENT_MODE= "0b0";
 parameter          RGB0_CURRENT= "0b000000";
 parameter          RGB1_CURRENT= "0b000000";
 parameter          RGB2_CURRENT= "0b000000";

//** Instantiate the  module **
SB_RGBA_DRV_CORE  #(.CURRENT_MODE(CURRENT_MODE), .RGB0_CURRENT(RGB0_CURRENT), .RGB1_CURRENT(RGB1_CURRENT), .RGB2_CURRENT(RGB2_CURRENT))
 inst_SB_RGBA_DRV    (
                      .RGB0PWM (RGB0PWM),
                      .RGB1PWM (RGB1PWM),
                      .RGB2PWM (RGB2PWM),
                      .CURREN (CURREN),
                      .RGBLEDEN (RGBLEDEN),

                      .RGB0 (RGB0),
                      .RGB1 (RGB1),
                      .RGB2 (RGB2));

`ifdef TIMINGCHECK
specify

   (RGB0PWM *> RGB0) = (1.0, 1.0);
   (RGB1PWM *> RGB1) = (1.0, 1.0);
   (RGB2PWM *> RGB2) = (1.0, 1.0);
   (RGBLEDEN *> RGB0) = (1.0, 1.0);
   (RGBLEDEN *> RGB1) = (1.0, 1.0);
   (RGBLEDEN *> RGB2) = (1.0, 1.0);

endspecify
`endif

endmodule

//--------------------------------------
// ----  SB_BARCODE_DRV ------ 
//--------------------------------------
`timescale 1ps/1ps
module SB_BARCODE_DRV   (
	CURREN,
	BARCODEEN,
	BARCODEPWM,
	BARCODE
);

parameter BARCODE_CURRENT = "0b0000";
parameter CURRENT_MODE = "0b0";

	input CURREN,	BARCODEEN, 	BARCODEPWM; 
	output 	BARCODE; 

 SB_BARCODE_DRV_CORE #(.BARCODE_CURRENT(BARCODE_CURRENT),.CURRENT_MODE(CURRENT_MODE))
inst
 (
	.CURREN(CURREN),
	.BARCODEEN(BARCODEEN),
	.BARCODEPWM(BARCODEPWM),
	.BARCODE(BARCODE)
);

`ifdef TIMINGCHECK
specify

   (BARCODEPWM *> BARCODE) = (1.0, 1.0);
   (BARCODEEN *> BARCODE) = (1.0, 1.0);
endspecify
`endif
endmodule

//--------------------------------------
// ----  SB_IR400_DRV ------ 
//--------------------------------------
`timescale 1ps/1ps
module SB_IR400_DRV   (
	CURREN,
	IRLEDEN,
	IRPWM,
	IRLED
);

parameter IR400_CURRENT = "0b00000000";
parameter CURRENT_MODE = "0b0";

	input CURREN,IRLEDEN,IRPWM;
	output 	IRLED; 

 SB_IR400_DRV_CORE #(.IR400_CURRENT(IR400_CURRENT),.CURRENT_MODE(CURRENT_MODE))
inst
 (
	.CURREN(CURREN),
	.IRLEDEN(IRLEDEN),
	.IRPWM(IRPWM),
	.IRLED(IRLED)
);
`ifdef TIMINGCHECK
specify

   (IRPWM *> IRLED) = (1.0, 1.0);
   (IRLEDEN *> IRLED) = (1.0, 1.0);
endspecify
`endif
endmodule
//--------------------------------------
// ----  SB_IR500_DRV ------ 
//--------------------------------------
`timescale 1ps/1ps
module SB_IR500_DRV   (
	IRLEDEN,
	IRPWM,
	CURREN,
	IRLED1,
	IRLED2
);

parameter IR500_CURRENT = "0b000000000000";
parameter CURRENT_MODE = "0b0";

	input IRLEDEN;
	input IRPWM;
	input CURREN;
	output IRLED1;
	output IRLED2;

 SB_IR500_DRV_CORE #(.IR500_CURRENT(IR500_CURRENT),.CURRENT_MODE(CURRENT_MODE))
inst
 (
	.CURREN(CURREN),
	.IRLEDEN(IRLEDEN),
	.IRPWM(IRPWM),
	.IRLED1(IRLED1),
	.IRLED2(IRLED2)
);
`ifdef TIMINGCHECK
specify

   (IRPWM *> IRLED1) = (1.0, 1.0);
   (IRPWM *> IRLED2) = (1.0, 1.0);
   (IRLEDEN *> IRLED1) = (1.0, 1.0);
   (IRLEDEN *> IRLED2) = (1.0, 1.0);
endspecify
`endif
endmodule

//--------------------------------------
// ----  SB_IR_IP ------ 
//--------------------------------------
`timescale 1ps/1ps
module SB_IR_IP(
// *** Input to UUT ***
 input            IRIN,
 input            ADRI3,
 input            ADRI2,
 input            ADRI1,
 input            ADRI0,
 input            CSI,
 input            DENI,
 input            EXE,
 input            LEARN,
 input            RST,
 input            WEI,
 input  		  CLKI,
// *** Outputs from UUT ***
 output            IROUT,
 output            BUSY,
 output            DRDY,
 output            ERR,
 output            RDATA0,
 output            RDATA1,
 output            RDATA2,
 output            RDATA3,
 output            RDATA4,
 output            RDATA5,
 output            RDATA6,
 output            RDATA7,


 input            WDATA0,
 input            WDATA1,
 input            WDATA2,
 input            WDATA3,
 input            WDATA4,
 input            WDATA5,
 input            WDATA6,
 input            WDATA7
 );

SB_IR_IP_CORE inst (
			 .CLKI(CLKI),
             .IRIN(IRIN),
             .ADRI3(ADRI3),
             .ADRI2(ADRI2),
             .ADRI1(ADRI1),
             .ADRI0(ADRI0),
             .CSI(CSI),
             .DENI(DENI),
             .EXE(EXE),
             .LEARN(LEARN),
             .RST(RST),
             .WEI(WEI),
             .IROUT(IROUT),
             .BUSY(BUSY),
             .DRDY(DRDY),
             .ERR(ERR),
             .RDATA0(RDATA0),
             .RDATA1(RDATA1),
             .RDATA2(RDATA2),
             .RDATA3(RDATA3),
             .RDATA4(RDATA4),
             .RDATA5(RDATA5),
             .RDATA6(RDATA6),
             .RDATA7(RDATA7),
             .WDATA0(WDATA0),
             .WDATA1(WDATA1),
             .WDATA2(WDATA2),
             .WDATA3(WDATA3),
             .WDATA4(WDATA4),
             .WDATA5(WDATA5),
             .WDATA6(WDATA6),
             .WDATA7(WDATA7)
);
`ifdef TIMINGCHECK
reg  NOTIFIER;
specify
	   $setuphold(posedge CLKI,posedge CSI,1.0,1.0, NOTIFIER);
       $setuphold( posedge CLKI,negedge CSI,1.0,1.0, NOTIFIER);
       $setuphold( posedge CLKI,posedge DENI,1.0,1.0, NOTIFIER);
       $setuphold( posedge CLKI,negedge DENI,1.0,1.0, NOTIFIER);
       $setuphold( posedge CLKI,posedge WEI,1.0,1.0, NOTIFIER);
       $setuphold( posedge CLKI,negedge WEI,1.0,1.0, NOTIFIER);
       $setuphold( posedge CLKI,posedge ADRI3,1.0,1.0, NOTIFIER);
       $setuphold( posedge CLKI,negedge ADRI3,1.0,1.0, NOTIFIER);
       $setuphold( posedge CLKI,posedge ADRI2,1.0,1.0, NOTIFIER);
       $setuphold( posedge CLKI,negedge ADRI2,1.0,1.0, NOTIFIER);
       $setuphold( posedge CLKI,posedge ADRI1,1.0,1.0, NOTIFIER);
       $setuphold( posedge CLKI,negedge ADRI1,1.0,1.0, NOTIFIER);
       $setuphold( posedge CLKI,posedge ADRI0,1.0,1.0, NOTIFIER);
       $setuphold( posedge CLKI,negedge ADRI0,1.0,1.0, NOTIFIER);
       $setuphold( posedge CLKI,posedge WDATA0,1.0,1.0, NOTIFIER);
       $setuphold( posedge CLKI,negedge WDATA0,1.0,1.0, NOTIFIER);
       $setuphold( posedge CLKI,posedge WDATA1,1.0,1.0, NOTIFIER);
       $setuphold( posedge CLKI,negedge WDATA1,1.0,1.0, NOTIFIER);
       $setuphold( posedge CLKI,posedge WDATA2,1.0,1.0, NOTIFIER);
       $setuphold( posedge CLKI,negedge WDATA2,1.0,1.0, NOTIFIER);
       $setuphold( posedge CLKI,posedge WDATA3,1.0,1.0, NOTIFIER);
       $setuphold( posedge CLKI,negedge WDATA3,1.0,1.0, NOTIFIER);
       $setuphold( posedge CLKI,posedge WDATA4,1.0,1.0, NOTIFIER);
       $setuphold( posedge CLKI,negedge WDATA4,1.0,1.0, NOTIFIER);
       $setuphold( posedge CLKI,posedge WDATA5,1.0,1.0, NOTIFIER);
       $setuphold( posedge CLKI,negedge WDATA5,1.0,1.0, NOTIFIER);
       $setuphold( posedge CLKI,posedge WDATA6,1.0,1.0, NOTIFIER);
       $setuphold( posedge CLKI,negedge WDATA6,1.0,1.0, NOTIFIER);
       $setuphold( posedge CLKI,posedge WDATA7,1.0,1.0, NOTIFIER);
       $setuphold( posedge CLKI,negedge WDATA7,1.0,1.0, NOTIFIER);
       $setuphold( posedge CLKI,posedge EXE,1.0,1.0, NOTIFIER);
       $setuphold( posedge CLKI,negedge EXE,1.0,1.0, NOTIFIER);
       $setuphold( posedge CLKI,posedge LEARN,1.0,1.0, NOTIFIER);
       $setuphold( posedge CLKI,negedge LEARN,1.0,1.0, NOTIFIER);
      (CLKI *> RDATA0)=(0.0,0.0);
      (CLKI *> RDATA1)=(0.0,0.0);
      (CLKI *> RDATA2)=(0.0,0.0);
      (CLKI *> RDATA3)=(0.0,0.0);
      (CLKI *> RDATA4)=(0.0,0.0);
      (CLKI *> RDATA5)=(0.0,0.0);
      (CLKI *> RDATA6)=(0.0,0.0);
      (CLKI *> RDATA7)=(0.0,0.0);
      (CLKI *> BUSY)=(0.0,0.0);
      (CLKI *> DRDY)=(0.0,0.0);
      (CLKI *> ERR)=(0.0,0.0);
      (CLKI *> IROUT)=(0.0,0.0);

endspecify
`endif
 endmodule
//--------------------------------------
// ----  SB_RGBA_DRV ------ 
//--------------------------------------
`timescale 1ps/1ps
module SB_I2C_FIFO (
input  CLKI,
input  CSI,
input  WEI,
input  STBI,
input  ADRI3,
input  ADRI2,
input  ADRI1,
input  ADRI0,
input  DATI0,
input  DATI1,
input  DATI2,
input  DATI3,
input  DATI4,
input  DATI5,
input  DATI6,
input  DATI7,
input  DATI8,
input  DATI9,
input  SCLI,
input  SDAI,
input  FIFORST,

output DATO0,
output DATO1,
output DATO2,
output DATO3,
output DATO4,
output DATO5,
output DATO6,
output DATO7,
output DATO8,
output DATO9,
output ACKO,
output I2CIRQ,
output I2CWKUP,
inout SCLO,
output SCLOE,
output SDAO,
output SDAOE,
output SRWO,
output	TXFIFOAEMPTY,
output	TXFIFOEMPTY,
output	TXFIFOFULL,
output	RXFIFOAFULL,
output	RXFIFOFULL,
output	RXFIFOEMPTY,
output MRDCMPL);


  parameter I2C_SLAVE_ADDR = "0b1111100001";
  //parameter BUS_ADDR74 = "0b0001";


wire master, slave;
assign (weak0, weak1) DATI0 =1'b0 ;
assign (weak0, weak1) DATI1 =1'b0 ;
assign (weak0, weak1) DATI2 =1'b0 ;
assign (weak0, weak1) DATI3 =1'b0 ;
assign (weak0, weak1) DATI4 =1'b0 ;
assign (weak0, weak1) DATI5 =1'b0 ;
assign (weak0, weak1) DATI6 =1'b0 ;
assign (weak0, weak1) DATI7 =1'b0 ;
assign (weak0, weak1) DATI8 =1'b0 ;
assign (weak0, weak1) DATI9 =1'b0 ;



SB_I2C_FIFO_CORE inst (
 	.CLKI(CLKI),
	.CSI(CSI),
 	.WEI(WEI),
 	.STBI(STBI),
 	.ADRI3(ADRI3),
 	.ADRI2(ADRI2),
 	.ADRI1(ADRI1),
 	.ADRI0(ADRI0),
	.DATI9(DATI9),
 	.DATI8(DATI8),
 	.DATI7(DATI7),
 	.DATI6(DATI6),
 	.DATI5(DATI5),
 	.DATI4(DATI4),
 	.DATI3(DATI3),
 	.DATI2(DATI2),
 	.DATI1(DATI1),
 	.DATI0(DATI0),
 	.SCLI(SCLI),
 	.SDAI(SDAI),
	.FIFORST(FIFORST),

	.DATO9(DATO9),
	.DATO8(DATO8),
	.DATO7(DATO7),
	.DATO6(DATO6),
	.DATO5(DATO5),
	.DATO4(DATO4),
	.DATO3(DATO3),
	.DATO2(DATO2),
	.DATO1(DATO1),
	.DATO0(DATO0),
	.ACKO(ACKO),
	.I2CIRQ(I2CIRQ),
	.I2CWKUP(I2CWKUP),
	.SCLO(SCLO),
	.SCLOE(SCLOE),
	.SDAO(SDAO),
	.SDAOE(SDAOE),
	.SRWO(SRWO),
  .TXFIFOAEMPTY(TXFIFOAEMPTY),
  .TXFIFOEMPTY(TXFIFOEMPTY),
  .TXFIFOFULL(TXFIFOFULL),
  .RXFIFOEMPTY(RXFIFOEMPTY),
  .RXFIFOAFULL(RXFIFOAFULL),
  .RXFIFOFULL(RXFIFOFULL),
	.MRDCMPL(MRDCMPL));
  defparam inst.I2C_SLAVE_ADDR = I2C_SLAVE_ADDR;
  //defparam inst.BUS_ADDR74 = BUS_ADDR74;

// initial begin
	// if (BUS_ADDR74!="0b0001" && BUS_ADDR74!="0b0011")
// $display ("ID:BUS_ADDR74: should be LLC=0b0001 or LRC=0b0011, otherwise there would be an error ");
// end

`ifdef TIMINGCHECK

reg NOTIFIER;
specify

   //(CLKI *> SCLO) = (1.0, 1.0);

   (CLKI *> TXFIFOAEMPTY) = (1.0, 1.0);
   (CLKI *> TXFIFOEMPTY) = (1.0, 1.0);
   (CLKI *> TXFIFOFULL) = (1.0, 1.0);
   (CLKI *> RXFIFOEMPTY) = (1.0, 1.0);
   (CLKI *> RXFIFOAFULL) = (1.0, 1.0);
   (CLKI *> RXFIFOFULL) = (1.0, 1.0);   
   (CLKI *> DATO0) = (1.0, 1.0);
   (CLKI *> DATO1) = (1.0, 1.0);
   (CLKI *> DATO2) = (1.0, 1.0);
   (CLKI *> DATO3) = (1.0, 1.0);
   (CLKI *> DATO4) = (1.0, 1.0);
   (CLKI *> DATO5) = (1.0, 1.0);
   (CLKI *> DATO6) = (1.0, 1.0);
   (CLKI *> DATO7) = (1.0, 1.0);
   (CLKI *> DATO8) = (1.0, 1.0);
   (CLKI *> DATO9) = (1.0, 1.0);
   (CLKI *> ACKO) = (1.0, 1.0);
   (CLKI *> SRWO) = (1.0, 1.0);
   (CLKI *> I2CIRQ) = (1.0, 1.0);
   (CLKI *> I2CWKUP) = (1.0, 1.0);
	(CLKI *> SCLO) = (1.0, 1.0);
	(CLKI *> SCLOE) = (1.0, 1.0);
    (SCLO *> SDAO) = (1.0, 1.0);
    (SCLO *> SDAOE) = (1.0, 1.0);
    (SCLI *> SDAO) = (1.0, 1.0);
    (SCLI *> SDAOE) = (1.0, 1.0);

   $setup(posedge WEI, posedge CLKI, 1.0);
   $setup(negedge WEI, posedge CLKI, 1.0);
   $hold(posedge CLKI, posedge WEI, 1.0);
   $hold(posedge CLKI, negedge WEI, 1.0);	 

   $setup(posedge STBI, posedge CLKI, 1.0);
   $setup(negedge STBI, posedge CLKI, 1.0);
   $hold(posedge CLKI, posedge STBI, 1.0);
   $hold(posedge CLKI, negedge STBI, 1.0);

   $setup(posedge CSI, posedge CLKI, 1.0);
   $setup(negedge CSI, posedge CLKI, 1.0);
   $hold(posedge CLKI, posedge CSI, 1.0);
   $hold(posedge CLKI, negedge CSI, 1.0);
   
   $setup(posedge FIFORST, posedge CLKI, 1.0);
   $setup(negedge FIFORST, posedge CLKI, 1.0);
   $hold(posedge CLKI, posedge FIFORST, 1.0);
   $hold(posedge CLKI, negedge FIFORST, 1.0);
   
   $setup(posedge SCLI, posedge CLKI, 1.0);
   $setup(negedge SCLI, posedge CLKI, 1.0);
   $hold(posedge CLKI, posedge SCLI, 1.0);
   $hold(posedge CLKI, negedge SCLI, 1.0); 
  
   $setup(posedge SDAI, posedge CLKI, 1.0);
   $setup(negedge SDAI, posedge CLKI, 1.0);
   $hold(posedge CLKI, posedge SDAI, 1.0);
   $hold(posedge CLKI, negedge SDAI, 1.0);
   
   $setup(posedge ADRI3, posedge CLKI, 1.0);
   $setup(negedge ADRI3, posedge CLKI, 1.0);
   $hold(posedge CLKI, posedge ADRI3, 1.0);
   $hold(posedge CLKI, negedge ADRI3, 1.0);

   $setup(posedge ADRI2, posedge CLKI, 1.0);
   $setup(negedge ADRI2, posedge CLKI, 1.0);
   $hold(posedge CLKI, posedge ADRI2, 1.0);
   $hold(posedge CLKI, negedge ADRI2, 1.0);

   $setup(posedge ADRI1, posedge CLKI, 1.0);
   $setup(negedge ADRI1, posedge CLKI, 1.0);
   $hold(posedge CLKI, posedge ADRI1, 1.0);
   $hold(posedge CLKI, negedge ADRI1, 1.0);

   $setup(posedge ADRI0, posedge CLKI, 1.0);
   $setup(negedge ADRI0, posedge CLKI, 1.0);
   $hold(posedge CLKI, posedge ADRI0, 1.0);
   $hold(posedge CLKI, negedge ADRI0, 1.0);

   
   $setup(posedge DATI9, posedge CLKI, 1.0);
   $setup(negedge DATI9, posedge CLKI, 1.0);
   $hold(posedge CLKI, posedge DATI9, 1.0);
   $hold(posedge CLKI, negedge DATI9, 1.0);
   
   
   $setup(posedge DATI8, posedge CLKI, 1.0);
   $setup(negedge DATI8, posedge CLKI, 1.0);
   $hold(posedge CLKI, posedge DATI8, 1.0);
   $hold(posedge CLKI, negedge DATI8, 1.0);
   
   $setup(posedge DATI7, posedge CLKI, 1.0);
   $setup(negedge DATI7, posedge CLKI, 1.0);
   $hold(posedge CLKI, posedge DATI7, 1.0);
   $hold(posedge CLKI, negedge DATI7, 1.0);

   $setup(posedge DATI6, posedge CLKI, 1.0);
   $setup(negedge DATI6, posedge CLKI, 1.0);
   $hold(posedge CLKI, posedge DATI6, 1.0);
   $hold(posedge CLKI, negedge DATI6, 1.0);

   $setup(posedge DATI5, posedge CLKI, 1.0);
   $setup(negedge DATI5, posedge CLKI, 1.0);
   $hold(posedge CLKI, posedge DATI5, 1.0);
   $hold(posedge CLKI, negedge DATI5, 1.0);

   $setup(posedge DATI4, posedge CLKI, 1.0);
   $setup(negedge DATI4, posedge CLKI, 1.0);
   $hold(posedge CLKI, posedge DATI4, 1.0);
   $hold(posedge CLKI, negedge DATI4, 1.0);

   $setup(posedge DATI3, posedge CLKI, 1.0);
   $setup(negedge DATI3, posedge CLKI, 1.0);
   $hold(posedge CLKI, posedge DATI3, 1.0);
   $hold(posedge CLKI, negedge DATI3, 1.0);

   $setup(posedge DATI2, posedge CLKI, 1.0);
   $setup(negedge DATI2, posedge CLKI, 1.0);
   $hold(posedge CLKI, posedge DATI2, 1.0);
   $hold(posedge CLKI, negedge DATI2, 1.0);

   $setup(posedge DATI1, posedge CLKI, 1.0);
   $setup(negedge DATI1, posedge CLKI, 1.0);
   $hold(posedge CLKI, posedge DATI1, 1.0);
   $hold(posedge CLKI, negedge DATI1, 1.0);

   $setup(posedge DATI0, posedge CLKI, 1.0);
   $setup(negedge DATI0, posedge CLKI, 1.0);
   $hold(posedge CLKI, posedge DATI0, 1.0);
   $hold(posedge CLKI, negedge DATI0, 1.0);

   $setuphold(posedge SCLO, posedge SDAI, 1.0, 1.0, NOTIFIER);
   $setuphold(posedge SCLO, negedge SDAI, 1.0, 1.0, NOTIFIER);

   $setuphold(posedge SCLI, posedge SDAI, 1.0, 1.0, NOTIFIER);
   $setuphold(posedge SCLI, negedge SDAI, 1.0, 1.0, NOTIFIER);

endspecify
`endif


endmodule


//-------------------------------------
// ----  SB_LEDDA_IP ------ 
//--------------------------------------
`timescale 1ps/1ps
module SB_LEDDA_IP ( LEDDCS,LEDDCLK,LEDDDAT7,LEDDDAT6,LEDDDAT5,LEDDDAT4,
	LEDDDAT3,LEDDDAT2,LEDDDAT1,LEDDDAT0,LEDDADDR3,LEDDADDR2,LEDDADDR1,
	LEDDADDR0,LEDDDEN,LEDDEXE,LEDDRST,PWMOUT0,PWMOUT1,PWMOUT2,LEDDON);	 
	
	input 	LEDDCS,LEDDCLK,LEDDDAT7,LEDDDAT6,LEDDDAT5,LEDDDAT4,LEDDDAT3,LEDDDAT2,
			LEDDDAT1,LEDDDAT0,LEDDADDR3,LEDDADDR2,LEDDADDR1,LEDDADDR0,LEDDDEN,LEDDEXE,LEDDRST; 
	output  PWMOUT0,PWMOUT1,PWMOUT2,LEDDON;
	
	wire LEDDCS, LEDDCLK,LEDDDAT7,LEDDDAT6,LEDDDAT5,LEDDDAT4,LEDDDAT3,LEDDDAT2, LEDDDAT1,LEDDDAT0,LEDDADDR3,LEDDADDR2,LEDDADDR1,LEDDADDR0,LEDDDEN,LEDDEXE,LEDDRST; 
	wire PWMOUT0,PWMOUT1,PWMOUT2,LEDDON;
	wire [7:0]  sb_ledd_dat={LEDDDAT7,LEDDDAT6,LEDDDAT5, LEDDDAT4,LEDDDAT3,LEDDDAT2,LEDDDAT1,LEDDDAT0};
	wire [3:0]	sb_ledd_adr={LEDDADDR3,LEDDADDR2,LEDDADDR1,LEDDADDR0};
	reg NOTIFIER;
	reg ledd_rst_async;
	initial
begin
   ledd_rst_async = 1'b1;
#100
   ledd_rst_async = 1'b0;
end
	ledd_ip  ledd_ip_inst
	(
	.pwm_out_r(PWMOUT0),
	.pwm_out_g(PWMOUT1), 
	.pwm_out_b(PWMOUT2), 
	.ledd_on(LEDDON),
	.ledd_rst_async(ledd_rst_async), 
	.ledd_clk(LEDDCLK), 
	.ledd_cs(LEDDCS), 
	.ledd_den(LEDDDEN), 
	.ledd_adr(sb_ledd_adr), 
	.ledd_dat(sb_ledd_dat),
    .ledd_exe(LEDDEXE)
   );
   
   `ifdef TIMINGCHECK
specify


	(LEDDCLK*>PWMOUT0) = (1.0, 1.0);
	(LEDDCLK*>PWMOUT1) = (1.0, 1.0);
	(LEDDCLK*>PWMOUT2) = (1.0, 1.0);
	(LEDDCLK*>LEDDON) = (1.0, 1.0);	 
   	$setup(posedge LEDDCS, posedge LEDDCLK,  1.0);  
	$setup(negedge LEDDCS, posedge LEDDCLK,  1.0); 
	$hold(posedge LEDDCLK, posedge LEDDCS,  1.0);
	$hold(posedge LEDDCLK, negedge LEDDCS,  1.0); 
	$setup(posedge LEDDDEN, posedge LEDDCLK,  1.0);  
	$setup(negedge LEDDDEN, posedge LEDDCLK,  1.0); 
	$hold(posedge LEDDCLK, posedge LEDDDEN,  1.0);
	$hold(posedge LEDDCLK, negedge LEDDDEN,  1.0);
	$setup(posedge LEDDEXE, posedge LEDDCLK,  1.0);  
	$setup(negedge LEDDEXE, posedge LEDDCLK,  1.0); 
	$hold(posedge LEDDCLK, posedge LEDDEXE,  1.0);
	$hold(posedge LEDDCLK, negedge LEDDEXE,  1.0);
	$setup(posedge LEDDADDR0, posedge LEDDCLK,  1.0);  
	$setup(negedge LEDDADDR0, posedge LEDDCLK,  1.0); 
	$hold(posedge LEDDCLK, posedge LEDDADDR0,  1.0);
	$hold(posedge LEDDCLK, negedge LEDDADDR0,  1.0);
	$setup(posedge LEDDADDR1, posedge LEDDCLK,  1.0);  
	$setup(negedge LEDDADDR1, posedge LEDDCLK,  1.0); 
	$hold(posedge LEDDCLK, posedge LEDDADDR1,  1.0);
	$hold(posedge LEDDCLK, negedge LEDDADDR1,  1.0);
	$setup(posedge LEDDADDR2, posedge LEDDCLK,  1.0);  
	$setup(negedge LEDDADDR2, posedge LEDDCLK,  1.0); 
	$hold(posedge LEDDCLK, posedge LEDDADDR2,  1.0);
	$hold(posedge LEDDCLK, negedge LEDDADDR2,  1.0);
	$setup(posedge LEDDADDR3, posedge LEDDCLK,  1.0);  
	$setup(negedge LEDDADDR3, posedge LEDDCLK,  1.0); 
	$hold(posedge LEDDCLK, posedge LEDDADDR3,  1.0);
	$hold(posedge LEDDCLK, negedge LEDDADDR3,  1.0);

	$setup(posedge LEDDDAT0, posedge LEDDCLK,  1.0);  
	$setup(negedge LEDDDAT0, posedge LEDDCLK,  1.0); 
	$hold(posedge LEDDCLK, posedge LEDDDAT0,  1.0);
	$hold(posedge LEDDCLK, negedge LEDDDAT0,  1.0);
	$setup(posedge LEDDDAT1, posedge LEDDCLK,  1.0);  
	$setup(negedge LEDDDAT1, posedge LEDDCLK,  1.0); 
	$hold(posedge LEDDCLK, posedge LEDDDAT1,  1.0);
	$hold(posedge LEDDCLK, negedge LEDDDAT1,  1.0);
	$setup(posedge LEDDDAT2, posedge LEDDCLK,  1.0);  
	$setup(negedge LEDDDAT2, posedge LEDDCLK,  1.0); 
	$hold(posedge LEDDCLK, posedge LEDDDAT2,  1.0);
	$hold(posedge LEDDCLK, negedge LEDDDAT2,  1.0);
	$setup(posedge LEDDDAT3, posedge LEDDCLK,  1.0);  
	$setup(negedge LEDDDAT3, posedge LEDDCLK,  1.0); 
	$hold(posedge LEDDCLK, posedge LEDDDAT3,  1.0);
	$hold(posedge LEDDCLK, negedge LEDDDAT3,  1.0);
	$setup(posedge LEDDDAT4, posedge LEDDCLK,  1.0);  
	$setup(negedge LEDDDAT4, posedge LEDDCLK,  1.0); 
	$hold(posedge LEDDCLK, posedge LEDDDAT4,  1.0);
	$hold(posedge LEDDCLK, negedge LEDDDAT4,  1.0);
	$setup(posedge LEDDDAT5, posedge LEDDCLK,  1.0);  
	$setup(negedge LEDDDAT5, posedge LEDDCLK,  1.0); 
	$hold(posedge LEDDCLK, posedge LEDDDAT5,  1.0);
	$hold(posedge LEDDCLK, negedge LEDDDAT5,  1.0);
	$setup(posedge LEDDDAT6, posedge LEDDCLK,  1.0);  
	$setup(negedge LEDDDAT6, posedge LEDDCLK,  1.0); 
	$hold(posedge LEDDCLK, posedge LEDDDAT6,  1.0);
	$hold(posedge LEDDCLK, negedge LEDDDAT6,  1.0);
	$setup(posedge LEDDDAT7, posedge LEDDCLK,  1.0);  
	$setup(negedge LEDDDAT7, posedge LEDDCLK,  1.0); 
	$hold(posedge LEDDCLK, posedge LEDDDAT7,  1.0);
	$hold(posedge LEDDCLK, negedge LEDDDAT7,  1.0);

		 endspecify
`endif

   
endmodule

//-------------------------------------
// ----  SB_RGB_IP ------ 
//--------------------------------------
`timescale 1ps/1ps
module  SB_RGB_IP ( 
CLK,RST,PARAMSOK,RGBCOLOR,BRIGHTNESS,BREATHRAMP,BLINKRATE,REDPWM,GREENPWM,BLUEPWM
); 
	input CLK; 
	input RST; 			
	input PARAMSOK; 
	input [3:0]  RGBCOLOR; 
	input [3:0] BRIGHTNESS; 
	input [3:0]BREATHRAMP; 
	input [3:0] BLINKRATE; 
	output REDPWM; 
	output GREENPWM; 
	output BLUEPWM;

LED_control RGBPWMinst (
       .clk27M(CLK),        
       .rst(RST),           
       .params_ok(PARAMSOK),     
       .RGB_color(RGBCOLOR),     
       .Brightness(BRIGHTNESS),    
       .BreatheRamp(BREATHRAMP),   
       .BlinkRate(BLINKRATE),     
       .red_pwm (REDPWM),       
       .grn_pwm(GREENPWM),       
       .blu_pwm(BLUEPWM)        
        );


endmodule 

//-------------------------------------
// ----  SB_SPRAM256KA ------ 
//--------------------------------------
`timescale 1ps / 1ps
module SB_SPRAM256KA(ADDRESS, DATAIN, MASKWREN,WREN,CHIPSELECT,CLOCK,STANDBY,SLEEP,POWEROFF,DATAOUT);
input [13:0] ADDRESS;
input [15:0] DATAIN;
input [3:0] MASKWREN;
input WREN,CHIPSELECT,CLOCK,STANDBY,SLEEP,POWEROFF;
output [15:0] DATAOUT;

wire [15:0]wem = {MASKWREN[3],MASKWREN[3],MASKWREN[3],MASKWREN[3],
					MASKWREN[2],MASKWREN[2],MASKWREN[2],MASKWREN[2],
					MASKWREN[1],MASKWREN[1],MASKWREN[1],MASKWREN[1],
					MASKWREN[0],MASKWREN[0],MASKWREN[0],MASKWREN[0]};

	
wire not_poweroff; 


assign (weak0, weak1) STANDBY 	=1'b0 ;
assign (weak0, weak1) SLEEP	=1'b0 ;
assign (weak0, weak1) POWEROFF 	=1'b1 ;			// Note: 1'b0-> POWEROFF, 1'b1 -> POWERON at wrapper level. 

assign not_poweroff = ~POWEROFF; 

sadslspk4s1p16384x16m16b4w1c0p1d0t0  spram256k_core_inst (
		.Q(DATAOUT),
		.ADR(ADDRESS),
		.D(DATAIN),
		.WEM(wem),
		.WE(WREN),
		.ME(CHIPSELECT),
		.CLK(CLOCK),
		.TEST1(),
		.RME(),
		.RM(),
		.LS(STANDBY),
		.DS(SLEEP),
		.SD(not_poweroff));	

`ifdef TIMINGCHECK
specify
	(CLOCK *> DATAOUT) = (1.0, 1.0);
	(SLEEP *> DATAOUT) = (1.0, 1.0);
   	$setup(posedge ADDRESS[0], posedge CLOCK,  1.0);  
	$setup(negedge ADDRESS[0], posedge CLOCK,  1.0); 
	$hold(posedge CLOCK, posedge ADDRESS[0],  1.0);
	$hold(posedge CLOCK, negedge ADDRESS[0],  1.0); 
   	$setup(posedge ADDRESS[1], posedge CLOCK,  1.0);  
	$setup(negedge ADDRESS[1], posedge CLOCK,  1.0); 
	$hold(posedge CLOCK, posedge ADDRESS[1],  1.0);
	$hold(posedge CLOCK, negedge ADDRESS[1],  1.0); 
   	$setup(posedge ADDRESS[2], posedge CLOCK,  1.0);  
	$setup(negedge ADDRESS[2], posedge CLOCK,  1.0); 
	$hold(posedge CLOCK, posedge ADDRESS[2],  1.0);
	$hold(posedge CLOCK, negedge ADDRESS[2],  1.0); 
   	$setup(posedge ADDRESS[3], posedge CLOCK,  1.0);  
	$setup(negedge ADDRESS[3], posedge CLOCK,  1.0); 
	$hold(posedge CLOCK, posedge ADDRESS[3],  1.0);
	$hold(posedge CLOCK, negedge ADDRESS[3],  1.0); 
   	$setup(posedge ADDRESS[4], posedge CLOCK,  1.0);  
	$setup(negedge ADDRESS[4], posedge CLOCK,  1.0); 
	$hold(posedge CLOCK, posedge ADDRESS[4],  1.0);
	$hold(posedge CLOCK, negedge ADDRESS[4],  1.0); 
   	$setup(posedge ADDRESS[5], posedge CLOCK,  1.0);  
	$setup(negedge ADDRESS[5], posedge CLOCK,  1.0); 
	$hold(posedge CLOCK, posedge ADDRESS[5],  1.0);
	$hold(posedge CLOCK, negedge ADDRESS[5],  1.0); 
   	$setup(posedge ADDRESS[6], posedge CLOCK,  1.0);  
	$setup(negedge ADDRESS[6], posedge CLOCK,  1.0); 
	$hold(posedge CLOCK, posedge ADDRESS[6],  1.0);
	$hold(posedge CLOCK, negedge ADDRESS[6],  1.0); 
   	$setup(posedge ADDRESS[7], posedge CLOCK,  1.0);  
	$setup(negedge ADDRESS[7], posedge CLOCK,  1.0); 
	$hold(posedge CLOCK, posedge ADDRESS[7],  1.0);
	$hold(posedge CLOCK, negedge ADDRESS[7],  1.0); 
   	$setup(posedge ADDRESS[8], posedge CLOCK,  1.0);  
	$setup(negedge ADDRESS[8], posedge CLOCK,  1.0); 
	$hold(posedge CLOCK, posedge ADDRESS[8],  1.0);
	$hold(posedge CLOCK, negedge ADDRESS[8],  1.0); 
   	$setup(posedge ADDRESS[9], posedge CLOCK,  1.0);  
	$setup(negedge ADDRESS[9], posedge CLOCK,  1.0); 
	$hold(posedge CLOCK, posedge ADDRESS[9],  1.0);
	$hold(posedge CLOCK, negedge ADDRESS[9],  1.0); 
   	$setup(posedge ADDRESS[10], posedge CLOCK,  1.0);  
	$setup(negedge ADDRESS[10], posedge CLOCK,  1.0); 
	$hold(posedge CLOCK, posedge ADDRESS[10],  1.0);
	$hold(posedge CLOCK, negedge ADDRESS[10],  1.0); 
   	$setup(posedge ADDRESS[11], posedge CLOCK,  1.0);  
	$setup(negedge ADDRESS[11], posedge CLOCK,  1.0); 
	$hold(posedge CLOCK, posedge ADDRESS[11],  1.0);
	$hold(posedge CLOCK, negedge ADDRESS[11],  1.0); 
   	$setup(posedge ADDRESS[12], posedge CLOCK,  1.0);  
	$setup(negedge ADDRESS[12], posedge CLOCK,  1.0); 
	$hold(posedge CLOCK, posedge ADDRESS[12],  1.0);
	$hold(posedge CLOCK, negedge ADDRESS[12],  1.0); 
   	$setup(posedge ADDRESS[13], posedge CLOCK,  1.0);  
	$setup(negedge ADDRESS[13], posedge CLOCK,  1.0); 
	$hold(posedge CLOCK, posedge ADDRESS[13],  1.0);
	$hold(posedge CLOCK, negedge ADDRESS[13],  1.0); 

	$setup(posedge DATAIN[0], posedge CLOCK,  1.0);  
	$setup(negedge DATAIN[0], posedge CLOCK,  1.0); 
	$hold(posedge CLOCK, posedge DATAIN[0],  1.0);
	$hold(posedge CLOCK, negedge DATAIN[0],  1.0); 
	$setup(posedge DATAIN[1], posedge CLOCK,  1.0);  
	$setup(negedge DATAIN[1], posedge CLOCK,  1.0); 
	$hold(posedge CLOCK, posedge DATAIN[1],  1.0);
	$hold(posedge CLOCK, negedge DATAIN[1],  1.0); 
	$setup(posedge DATAIN[2], posedge CLOCK,  1.0);  
	$setup(negedge DATAIN[2], posedge CLOCK,  1.0); 
	$hold(posedge CLOCK, posedge DATAIN[2],  1.0);
	$hold(posedge CLOCK, negedge DATAIN[2],  1.0); 
	$setup(posedge DATAIN[3], posedge CLOCK,  1.0);  
	$setup(negedge DATAIN[3], posedge CLOCK,  1.0); 
	$hold(posedge CLOCK, posedge DATAIN[3],  1.0);
	$hold(posedge CLOCK, negedge DATAIN[3],  1.0); 
	$setup(posedge DATAIN[4], posedge CLOCK,  1.0);  
	$setup(negedge DATAIN[4], posedge CLOCK,  1.0); 
	$hold(posedge CLOCK, posedge DATAIN[4],  1.0);
	$hold(posedge CLOCK, negedge DATAIN[4],  1.0); 
	$setup(posedge DATAIN[5], posedge CLOCK,  1.0);  
	$setup(negedge DATAIN[5], posedge CLOCK,  1.0); 
	$hold(posedge CLOCK, posedge DATAIN[5],  1.0);
	$hold(posedge CLOCK, negedge DATAIN[5],  1.0); 
	$setup(posedge DATAIN[6], posedge CLOCK,  1.0);  
	$setup(negedge DATAIN[6], posedge CLOCK,  1.0); 
	$hold(posedge CLOCK, posedge DATAIN[6],  1.0);
	$hold(posedge CLOCK, negedge DATAIN[6],  1.0); 
	$setup(posedge DATAIN[7], posedge CLOCK,  1.0);  
	$setup(negedge DATAIN[7], posedge CLOCK,  1.0); 
	$hold(posedge CLOCK, posedge DATAIN[7],  1.0);
	$hold(posedge CLOCK, negedge DATAIN[7],  1.0); 
	$setup(posedge DATAIN[8], posedge CLOCK,  1.0);  
	$setup(negedge DATAIN[8], posedge CLOCK,  1.0); 
	$hold(posedge CLOCK, posedge DATAIN[8],  1.0);
	$hold(posedge CLOCK, negedge DATAIN[8],  1.0); 
	$setup(posedge DATAIN[9], posedge CLOCK,  1.0);  
	$setup(negedge DATAIN[9], posedge CLOCK,  1.0); 
	$hold(posedge CLOCK, posedge DATAIN[9],  1.0);
	$hold(posedge CLOCK, negedge DATAIN[9],  1.0); 
	$setup(posedge DATAIN[10], posedge CLOCK,  1.0);  
	$setup(negedge DATAIN[10], posedge CLOCK,  1.0); 
	$hold(posedge CLOCK, posedge DATAIN[10],  1.0);
	$hold(posedge CLOCK, negedge DATAIN[10],  1.0); 
	$setup(posedge DATAIN[11], posedge CLOCK,  1.0);  
	$setup(negedge DATAIN[11], posedge CLOCK,  1.0); 
	$hold(posedge CLOCK, posedge DATAIN[11],  1.0);
	$hold(posedge CLOCK, negedge DATAIN[11],  1.0); 
	$setup(posedge DATAIN[12], posedge CLOCK,  1.0);  
	$setup(negedge DATAIN[12], posedge CLOCK,  1.0); 
	$hold(posedge CLOCK, posedge DATAIN[12],  1.0);
	$hold(posedge CLOCK, negedge DATAIN[12],  1.0); 
	$setup(posedge DATAIN[13], posedge CLOCK,  1.0);  
	$setup(negedge DATAIN[13], posedge CLOCK,  1.0); 
	$hold(posedge CLOCK, posedge DATAIN[13],  1.0);
	$hold(posedge CLOCK, negedge DATAIN[13],  1.0); 
	$setup(posedge DATAIN[14], posedge CLOCK,  1.0);  
	$setup(negedge DATAIN[14], posedge CLOCK,  1.0); 
	$hold(posedge CLOCK, posedge DATAIN[14],  1.0);
	$hold(posedge CLOCK, negedge DATAIN[14],  1.0); 
	$setup(posedge DATAIN[15], posedge CLOCK,  1.0);  
	$setup(negedge DATAIN[15], posedge CLOCK,  1.0); 
	$hold(posedge CLOCK, posedge DATAIN[15],  1.0);
	$hold(posedge CLOCK, negedge DATAIN[15],  1.0); 

	$setup(posedge MASKWREN[0], posedge CLOCK,  1.0);  
	$setup(negedge MASKWREN[0], posedge CLOCK,  1.0); 
	$hold(posedge CLOCK, posedge MASKWREN[0],  1.0);
	$hold(posedge CLOCK, negedge MASKWREN[0],  1.0); 
	$setup(posedge MASKWREN[1], posedge CLOCK,  1.0);  
	$setup(negedge MASKWREN[1], posedge CLOCK,  1.0); 
	$hold(posedge CLOCK, posedge MASKWREN[1],  1.0);
	$hold(posedge CLOCK, negedge MASKWREN[1],  1.0); 
	$setup(posedge MASKWREN[2], posedge CLOCK,  1.0);  
	$setup(negedge MASKWREN[2], posedge CLOCK,  1.0); 
	$hold(posedge CLOCK, posedge MASKWREN[2],  1.0);
	$hold(posedge CLOCK, negedge MASKWREN[2],  1.0); 
	$setup(posedge MASKWREN[3], posedge CLOCK,  1.0);  
	$setup(negedge MASKWREN[3], posedge CLOCK,  1.0); 
	$hold(posedge CLOCK, posedge MASKWREN[3],  1.0);
	$hold(posedge CLOCK, negedge MASKWREN[3],  1.0); 

	$setup(posedge WREN, posedge CLOCK,  1.0);  
	$setup(negedge WREN, posedge CLOCK,  1.0); 
	$hold(posedge CLOCK, posedge WREN,  1.0);
	$hold(posedge CLOCK, negedge WREN,  1.0); 
	$setup(posedge CHIPSELECT, posedge CLOCK,  1.0);  
	$setup(negedge CHIPSELECT, posedge CLOCK,  1.0); 
	$hold(posedge CLOCK, posedge CHIPSELECT,  1.0);
	$hold(posedge CLOCK, negedge CHIPSELECT,  1.0);
	$setup(posedge STANDBY, posedge CLOCK,  1.0);  
	$setup(negedge STANDBY, posedge CLOCK,  1.0); 
	$hold(posedge CLOCK, posedge STANDBY,  1.0);
	$hold(posedge CLOCK, negedge STANDBY,  1.0);
	$setup(posedge SLEEP, posedge CLOCK,  1.0);  
	$setup(negedge SLEEP, posedge CLOCK,  1.0); 
	$hold(posedge CLOCK, posedge SLEEP,  1.0);
	$hold(posedge CLOCK, negedge SLEEP,  1.0);

endspecify
`endif

endmodule

//--------------------------------------------------------------//
//--------   SB_IO_I3C  ---------------------------------------// 
//-------------------------------------------------------------//


`timescale 10ps/1ps

module SB_IO_I3C (
	PACKAGE_PIN, 
	LATCH_INPUT_VALUE, 
	CLOCK_ENABLE, 
	INPUT_CLK, 
	OUTPUT_CLK, 
	OUTPUT_ENABLE, 
	D_OUT_1, 
	D_OUT_0, 
	D_IN_1, 
	D_IN_0 , 
	PU_ENB, 
	WEAK_PU_ENB
 );

parameter PIN_TYPE     = 6'b000000;	 
parameter PULLUP       = 1'b0;    	// By default PULL Up=0. Set  1'b1 to enable 3p3k/6p8k/10k resistors controlled by PU_ENB signal.           
parameter WEAK_PULLUP  = 1'b0;          // By default WEAK Pull Up=0. Set 1'b1 to enable 100K weak pullup resistor controlled by WEAK_PU_ENB signal.     
parameter NEG_TRIGGER  = 1'b0;            
parameter IO_STANDARD  = "SB_LVCMOS";     			 

input D_OUT_1;  			// Input output 1
input D_OUT_0;  			// Input output 0
input CLOCK_ENABLE;    			// Clock enables in/out clocks

output D_IN_1;    			// Output input 1
output D_IN_0;    			// Output input 0

input OUTPUT_ENABLE;   			// Ouput-Enable 
input LATCH_INPUT_VALUE;    		// Input control
input INPUT_CLK;   			// Input clock
input OUTPUT_CLK;  			// Output clock
inout PACKAGE_PIN; 			// User's package pin - 'PAD' output.

input PU_ENB; 				// Active low pullup resistor enable/disable signal.  
input WEAK_PU_ENB;			// Active low weak pullup resistor enable/disable signal.  


//------------- Main Body of verilog ----------------------------------------------------
wire inclk_, outclk_;
wire inclk, outclk;
reg INCLKE_sync, OUTCLKE_sync; 

assign (weak0, weak1) CLOCK_ENABLE =1'b1 ;
assign inclk_ = (INPUT_CLK ^ NEG_TRIGGER); 	// change the input clock phase
assign outclk_ = (OUTPUT_CLK ^ NEG_TRIGGER);	 // change the output clock phase

//////// CLKEN sync ///////
always@(inclk_ or CLOCK_ENABLE)
begin 
    if(~inclk_)
	INCLKE_sync = CLOCK_ENABLE; 
end

always@(outclk_ or CLOCK_ENABLE)
begin 
   if(~outclk_) 	
	OUTCLKE_sync = CLOCK_ENABLE; 
end

assign inclk = (inclk_ & INCLKE_sync);
assign outclk = (outclk_ & OUTCLKE_sync);

wire bs_en;   //Boundary scan enable
wire shift;   //Boundary scan shift
wire tclk;    //Boundary scan clock
wire update;  //Boundary scan update
wire sdi;     //Boundary scan serial data in
wire mode;    //Boundary scan mode
wire hiz_b;   //Boundary scan tristate control
wire sdo;     //Boundary scan serial data out


assign  bs_en = 1'b0;	//Boundary scan enable
assign  shift = 1'b0;	//Boundary scan shift
assign  tclk = 1'b0;	//Boundary scan clock
assign  update = 1'b0;	//Boundary scan update
assign  sdi = 1'b0;	//Boundary scan serial data in
assign  mode = 1'b0;	//Boundary scan mode
assign  hiz_b = 1'b1;	//Boundary scan Tristate control
  
wire padoen, padout, padin;
assign PACKAGE_PIN = (~padoen) ? padout : 1'bz;
assign padin = PACKAGE_PIN ;



wire hold, oepin;							  // The required package pin type must be set when io_macro is instantiated.
assign hold = LATCH_INPUT_VALUE;
assign oepin = OUTPUT_ENABLE;
 
 preio_physical preiophysical_i (	//original names unchanged
 	.hold(hold),
	.rstio(1'b0),			//Disabled as this is power on only.
	.bs_en(bs_en),
	.shift(shift),
	.tclk(tclk),
	.inclk(inclk),
	.outclk(outclk),
	.update(update),
	.oepin(oepin),
	.sdi(sdi),
	.mode(mode),
	.hiz_b(hiz_b),
	.sdo(sdo),
	.dout1(D_IN_1),
	.dout0(D_IN_0),
	.ddr1(D_OUT_1),
	.ddr0(D_OUT_0),
	.padin(padin),
	.padout(padout),
	.padoen(padoen),
	.cbit(PIN_TYPE)
	);

`ifdef TIMINGCHECK
specify

   (PACKAGE_PIN *> D_IN_0) = (1.0, 1.0);
   (PACKAGE_PIN *> D_IN_1) = (1.0, 1.0);
   (INPUT_CLK *> D_IN_0) = (1.0, 1.0);
   (INPUT_CLK *> D_IN_1) = (1.0, 1.0);
   (D_OUT_0 *> PACKAGE_PIN) = (1.0, 1.0);
   (D_OUT_1 *> PACKAGE_PIN) = (1.0, 1.0);
   (OUTPUT_ENABLE *> PACKAGE_PIN) = (1.0, 1.0);
   (INPUT_CLK *> PACKAGE_PIN) = (1.0, 1.0);
   (OUTPUT_CLK *> PACKAGE_PIN) = (1.0, 1.0);
   (LATCH_INPUT_VALUE *> D_IN_0) = (1.0, 1.0);
   (LATCH_INPUT_VALUE *> D_IN_1) = (1.0, 1.0);

   $setup(posedge CLOCK_ENABLE, posedge INPUT_CLK, 1.0);
   $setup(negedge CLOCK_ENABLE, posedge INPUT_CLK, 1.0);
   $hold(posedge INPUT_CLK, posedge CLOCK_ENABLE, 1.0);
   $hold(posedge INPUT_CLK, negedge CLOCK_ENABLE, 1.0);
   $setup(posedge PACKAGE_PIN, posedge INPUT_CLK, 1.0);
   $setup(negedge PACKAGE_PIN, posedge INPUT_CLK, 1.0);
   $hold(posedge INPUT_CLK, posedge PACKAGE_PIN, 1.0);
   $hold(posedge INPUT_CLK, negedge PACKAGE_PIN, 1.0);
   $setup(posedge PACKAGE_PIN, negedge INPUT_CLK, 1.0);
   $setup(negedge PACKAGE_PIN, negedge INPUT_CLK, 1.0);
   $hold(negedge INPUT_CLK, posedge PACKAGE_PIN, 1.0);
   $hold(negedge INPUT_CLK, negedge PACKAGE_PIN, 1.0);
   $setup(posedge CLOCK_ENABLE, posedge OUTPUT_CLK, 1.0);
   $setup(negedge CLOCK_ENABLE, posedge OUTPUT_CLK, 1.0);
   $hold(posedge OUTPUT_CLK, posedge CLOCK_ENABLE, 1.0);
   $hold(posedge OUTPUT_CLK, negedge CLOCK_ENABLE, 1.0);
   $setup(posedge PACKAGE_PIN, posedge OUTPUT_CLK, 1.0);
   $setup(negedge PACKAGE_PIN, posedge OUTPUT_CLK, 1.0);
   $hold(posedge OUTPUT_CLK, posedge PACKAGE_PIN, 1.0);
   $hold(posedge OUTPUT_CLK, negedge PACKAGE_PIN, 1.0);
   $setup(posedge D_OUT_0, posedge OUTPUT_CLK, 1.0);
   $setup(negedge D_OUT_0, posedge OUTPUT_CLK, 1.0);
   $hold(posedge OUTPUT_CLK, posedge D_OUT_0, 1.0);
   $hold(posedge OUTPUT_CLK, negedge D_OUT_0, 1.0);
   $setup(posedge D_OUT_1, posedge OUTPUT_CLK, 1.0);
   $setup(negedge D_OUT_1, posedge OUTPUT_CLK, 1.0);
   $hold(posedge OUTPUT_CLK, posedge D_OUT_1, 1.0);
   $hold(posedge OUTPUT_CLK, negedge D_OUT_1, 1.0);
   $setup(posedge D_OUT_1, negedge OUTPUT_CLK, 1.0);
   $setup(negedge D_OUT_1, negedge OUTPUT_CLK, 1.0);
   $hold(negedge OUTPUT_CLK, posedge D_OUT_1, 1.0);
   $hold(negedge OUTPUT_CLK, negedge D_OUT_1, 1.0);
   $setup(posedge D_OUT_0, posedge OUTPUT_CLK, 1.0);
   $setup(negedge D_OUT_0, posedge OUTPUT_CLK, 1.0);
   $hold(posedge OUTPUT_CLK, posedge D_OUT_0, 1.0);
   $hold(posedge OUTPUT_CLK, negedge D_OUT_0, 1.0);
   $setup(posedge OUTPUT_ENABLE, posedge OUTPUT_CLK, 1.0);
   $setup(negedge OUTPUT_ENABLE, posedge OUTPUT_CLK, 1.0);
   $hold(posedge OUTPUT_CLK, posedge OUTPUT_ENABLE, 1.0);
   $hold(posedge OUTPUT_CLK, negedge OUTPUT_ENABLE, 1.0);

endspecify
`endif

endmodule

//--------------------------------------------------------------//
//--------   SB_FILTER_50NS-------------------------------------// 
//-------------------------------------------------------------//
//------ Glitch Filter with 50Ns Delay -----------------------// 

module SB_FILTER_50NS ( 
			FILTERIN,	
			FILTEROUT 
			); 

input FILTERIN; 
output FILTEROUT; 


assign FILTEROUT=FILTERIN; 


`ifdef TIMINGCHECK
specify 

  (FILTERIN => FILTEROUT) = (1.0,1.0); 

endspecify
`endif

endmodule




// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.10.0.111.2
// Netlist written on Wed Jul 11 11:47:38 2018
//
// Verilog Description of module aes
//

module aes (clk, reset_n, cs, we, address, write_data, read_data) /* synthesis syn_module_defined=1 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(39[8:11])
    input clk;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(41[33:36])
    input reset_n;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(42[33:40])
    input cs;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(45[33:35])
    input we;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(46[33:35])
    input [7:0]address;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(49[33:40])
    input [31:0]write_data;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(50[33:43])
    output [31:0]read_data;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(51[33:42])
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(41[33:36])
    
    wire GND_net, VCC_net, result_valid_new, reset_n_c, cs_c, we_c, 
        address_c_7, address_c_6, address_c_5, address_c_4, address_c_3, 
        address_c_2, address_c_1, address_c_0, write_data_c_31, write_data_c_30, 
        write_data_c_29, write_data_c_28, write_data_c_27, write_data_c_26, 
        write_data_c_25, write_data_c_24, write_data_c_23, write_data_c_22, 
        write_data_c_21, write_data_c_20, write_data_c_19, write_data_c_18, 
        write_data_c_17, write_data_c_16, write_data_c_15, write_data_c_14, 
        write_data_c_13, write_data_c_12, write_data_c_11, write_data_c_10, 
        write_data_c_9, write_data_c_8, write_data_c_7, write_data_c_6, 
        write_data_c_5, write_data_c_4, write_data_c_3, write_data_c_2, 
        write_data_c_1, write_data_c_0, read_data_c_31, read_data_c_30, 
        read_data_c_29, read_data_c_28, read_data_c_27, read_data_c_26, 
        read_data_c_25, read_data_c_24, read_data_c_23, read_data_c_22, 
        read_data_c_21, read_data_c_20, read_data_c_19, read_data_c_18, 
        read_data_c_17, read_data_c_16, read_data_c_15, read_data_c_14, 
        read_data_c_13, read_data_c_12, read_data_c_11, read_data_c_10, 
        read_data_c_9, read_data_c_8, read_data_c_7, read_data_c_6, 
        read_data_c_5, read_data_c_4, read_data_c_3, read_data_c_2, 
        read_data_c_1, read_data_c_0, encdec_reg, config_we;
    wire [31:0]\block_reg[0] ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(100[16:25])
    wire [31:0]\block_reg[1] ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(100[16:25])
    wire [31:0]\block_reg[2] ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(100[16:25])
    wire [31:0]\block_reg[3] ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(100[16:25])
    wire [31:0]\key_reg[0] ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(103[16:23])
    wire [31:0]\key_reg[1] ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(103[16:23])
    wire [31:0]\key_reg[2] ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(103[16:23])
    wire [31:0]\key_reg[3] ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(103[16:23])
    wire [31:0]\key_reg[4] ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(103[16:23])
    wire [31:0]\key_reg[5] ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(103[16:23])
    wire [31:0]\key_reg[6] ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(103[16:23])
    wire [31:0]\key_reg[7] ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(103[16:23])
    wire [127:0]result_reg;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(106[17:27])
    
    wire valid_reg, ready_reg, core_ready;
    wire [127:0]core_result;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(123[18:29])
    
    wire core_valid, n17169, n17104, n17109, n16989, n17044, n17049, 
        n16984, n16864, n16869, n16804, n16809, n16744, n16749, 
        n16684, n16689, n1504, init_state, ready_we;
    wire [1:0]aes_core_ctrl_reg;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(71[15:32])
    
    wire result_valid_we;
    wire [3:0]dec_round_nr;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(99[18:30])
    wire [31:0]muxed_sboxw;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(109[18:29])
    wire [31:0]new_sboxw;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(110[18:27])
    wire [1:0]aes_core_ctrl_new_1__N_858;
    wire [3:0]round_ctr_new;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(201[17:30])
    
    wire round_ctr_we, n16624, n16629, dec_ctrl_we;
    wire [31:0]tmp_sboxw;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(228[17:26])
    wire [31:0]new_sboxw_adj_9440;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(229[17:26])
    
    wire n16564, n16569, n16504, n16509, n16444, n16449, n34046, 
        n34043, n34040, n34037, n34034, n34031, n34028, n34025, 
        n34022, n34019, n34016, n34013, n34010, n34007, n34004, 
        n34001, n33998, n33995, n33992, n33989, n33986, n28832, 
        dec_ctrl_new_2__N_2032, clk_c_enable_2540, clk_c_enable_2508, 
        clk_c_enable_2476, clk_c_enable_387, clk_c_enable_355, clk_c_enable_323, 
        clk_c_enable_291, clk_c_enable_259, clk_c_enable_227, n16384, 
        n28824, n16389, round_ctr_we_adj_9437, n16324, n16329, n28846, 
        n28841, n28831, n28830, n16264, n16269, n16204, n16209, 
        n16144, n16149, clk_c_enable_195, n16084, n33861, n33860, 
        n33858, n33857, n33850, n16089, enc_ctrl_new_2__N_1045, n16024, 
        n16029, n15964, n15969, n15904, n15909;
    wire [3:0]\key_mem_ctrl.num_rounds ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(366[19:29])
    
    wire n10461, n15844, n15849, n15784, n15789, n15724, n15729, 
        n15664, n15669, n15604, n15609, n15544, n15549, n15484, 
        n15489, n15424, n15429, n15362, n15316, n28845, n33954, 
        n33953, n152, n14930, n14934, n14939, n149, n37, n33, 
        n17164, n17224, n17229;
    wire [127:0]prev_key1_new_127__N_4787;
    wire [2:0]key_mem_ctrl_new_2__N_4928;
    
    wire clk_c_enable_2444, clk_c_enable_163, n16924, n16929, n13203, 
        n13202, n1, n33950, n33949, n33948, n33947, n33946, n33942, 
        n33941, n33940, n33939, n8904, n33956, n25954, n20756, 
        n33915, n33913, n33910, n33909, n34048, n34047, n34045, 
        n34044, n34042, n34041, n34039, n34038, n34036, n34035, 
        n34033, n34032, n34030, n34029, n34027, n34026, n34024, 
        n34023, n34021, n34020, n34018, n34017, n34015, n34014, 
        n34012, n34011, n34009, n34008, n34006, n34005, n34003, 
        n34002, n34000, n33999, n33997, n33996, n33994, n35835, 
        n33993, n33991, n33990, n33988, n33987, n33985, n33984, 
        n33983, n33981, n33980, n33978, n33977, n33975, n33974, 
        n33972, n33971, n33969, n33968, n33966, n33965, n33963, 
        n33962, n33960, n33959, n33957;
    
    VHI i30299 (.Z(VCC_net));
    FD1S3AX result_reg_i0 (.D(core_result[0]), .CK(clk_c), .Q(result_reg[0]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i0.GSR = "ENABLED";
    FD1S3AX valid_reg_108 (.D(core_valid), .CK(clk_c), .Q(valid_reg));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam valid_reg_108.GSR = "ENABLED";
    FD1S3AX ready_reg_109 (.D(core_ready), .CK(clk_c), .Q(ready_reg));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam ready_reg_109.GSR = "ENABLED";
    FD1P3AX key_reg_7___i1 (.D(write_data_c_0), .SP(clk_c_enable_163), .CK(clk_c), 
            .Q(\key_reg[7] [0]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i1.GSR = "ENABLED";
    FD1S3AX result_reg_i26 (.D(core_result[26]), .CK(clk_c), .Q(result_reg[26]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i26.GSR = "ENABLED";
    FD1S3AX result_reg_i25 (.D(core_result[25]), .CK(clk_c), .Q(result_reg[25]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i25.GSR = "ENABLED";
    FD1S3AX result_reg_i24 (.D(core_result[24]), .CK(clk_c), .Q(result_reg[24]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i24.GSR = "ENABLED";
    FD1S3AX result_reg_i23 (.D(core_result[23]), .CK(clk_c), .Q(result_reg[23]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i23.GSR = "ENABLED";
    FD1S3AX result_reg_i22 (.D(core_result[22]), .CK(clk_c), .Q(result_reg[22]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i22.GSR = "ENABLED";
    FD1S3AX result_reg_i21 (.D(core_result[21]), .CK(clk_c), .Q(result_reg[21]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i21.GSR = "ENABLED";
    FD1S3AX result_reg_i20 (.D(core_result[20]), .CK(clk_c), .Q(result_reg[20]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i20.GSR = "ENABLED";
    FD1S3AX result_reg_i19 (.D(core_result[19]), .CK(clk_c), .Q(result_reg[19]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i19.GSR = "ENABLED";
    FD1S3AX result_reg_i18 (.D(core_result[18]), .CK(clk_c), .Q(result_reg[18]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i18.GSR = "ENABLED";
    FD1S3AX result_reg_i17 (.D(core_result[17]), .CK(clk_c), .Q(result_reg[17]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i17.GSR = "ENABLED";
    FD1S3AX result_reg_i16 (.D(core_result[16]), .CK(clk_c), .Q(result_reg[16]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i16.GSR = "ENABLED";
    FD1S3AX result_reg_i15 (.D(core_result[15]), .CK(clk_c), .Q(result_reg[15]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i15.GSR = "ENABLED";
    FD1S3AX result_reg_i14 (.D(core_result[14]), .CK(clk_c), .Q(result_reg[14]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i14.GSR = "ENABLED";
    FD1S3AX result_reg_i13 (.D(core_result[13]), .CK(clk_c), .Q(result_reg[13]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i13.GSR = "ENABLED";
    FD1S3AX result_reg_i12 (.D(core_result[12]), .CK(clk_c), .Q(result_reg[12]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i12.GSR = "ENABLED";
    FD1S3AX result_reg_i11 (.D(core_result[11]), .CK(clk_c), .Q(result_reg[11]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i11.GSR = "ENABLED";
    FD1S3AX result_reg_i10 (.D(core_result[10]), .CK(clk_c), .Q(result_reg[10]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i10.GSR = "ENABLED";
    FD1S3AX result_reg_i9 (.D(core_result[9]), .CK(clk_c), .Q(result_reg[9]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i9.GSR = "ENABLED";
    FD1S3AX result_reg_i8 (.D(core_result[8]), .CK(clk_c), .Q(result_reg[8]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i8.GSR = "ENABLED";
    FD1S3AX result_reg_i7 (.D(core_result[7]), .CK(clk_c), .Q(result_reg[7]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i7.GSR = "ENABLED";
    FD1S3AX result_reg_i6 (.D(core_result[6]), .CK(clk_c), .Q(result_reg[6]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i6.GSR = "ENABLED";
    FD1S3AX result_reg_i5 (.D(core_result[5]), .CK(clk_c), .Q(result_reg[5]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i5.GSR = "ENABLED";
    FD1S3AX result_reg_i4 (.D(core_result[4]), .CK(clk_c), .Q(result_reg[4]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i4.GSR = "ENABLED";
    FD1S3AX result_reg_i3 (.D(core_result[3]), .CK(clk_c), .Q(result_reg[3]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i3.GSR = "ENABLED";
    FD1S3AX result_reg_i2 (.D(core_result[2]), .CK(clk_c), .Q(result_reg[2]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i2.GSR = "ENABLED";
    FD1S3AX result_reg_i1 (.D(core_result[1]), .CK(clk_c), .Q(result_reg[1]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i1.GSR = "ENABLED";
    LUT4 n30951_bdd_4_lut_4_lut_then_4_lut (.A(n8904), .B(address_c_0), 
         .C(result_reg[11]), .D(result_reg[43]), .Z(n33957)) /* synthesis lut_function=(A (B (C)+!B (D))) */ ;
    defparam n30951_bdd_4_lut_4_lut_then_4_lut.init = 16'ha280;
    LUT4 n30951_bdd_4_lut_4_lut_else_4_lut (.A(n8904), .B(result_reg[75]), 
         .C(result_reg[107]), .D(address_c_0), .Z(n33956)) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam n30951_bdd_4_lut_4_lut_else_4_lut.init = 16'h88a0;
    PFUMX i29078 (.BLUT(n34043), .ALUT(n34044), .C0(address_c_1), .Z(n34045));
    PFUMX i29076 (.BLUT(n34040), .ALUT(n34041), .C0(address_c_0), .Z(n34042));
    LUT4 n30936_bdd_4_lut_4_lut_then_4_lut (.A(n8904), .B(address_c_0), 
         .C(result_reg[6]), .D(result_reg[38]), .Z(n33960)) /* synthesis lut_function=(A (B (C)+!B (D))) */ ;
    defparam n30936_bdd_4_lut_4_lut_then_4_lut.init = 16'ha280;
    PFUMX i29074 (.BLUT(n34037), .ALUT(n34038), .C0(address_c_0), .Z(n34039));
    LUT4 n30936_bdd_4_lut_4_lut_else_4_lut (.A(n8904), .B(result_reg[70]), 
         .C(result_reg[102]), .D(address_c_0), .Z(n33959)) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam n30936_bdd_4_lut_4_lut_else_4_lut.init = 16'h88a0;
    LUT4 i2_3_lut (.A(address_c_7), .B(address_c_5), .C(address_c_6), 
         .Z(n15362)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(49[33:40])
    defparam i2_3_lut.init = 16'hfefe;
    PFUMX i29072 (.BLUT(n34034), .ALUT(n34035), .C0(address_c_0), .Z(n34036));
    PFUMX i29070 (.BLUT(n34031), .ALUT(n34032), .C0(address_c_0), .Z(n34033));
    PFUMX i29068 (.BLUT(n34028), .ALUT(n34029), .C0(address_c_0), .Z(n34030));
    LUT4 n30987_bdd_4_lut_4_lut_then_4_lut (.A(n8904), .B(address_c_0), 
         .C(result_reg[23]), .D(result_reg[55]), .Z(n33963)) /* synthesis lut_function=(A (B (C)+!B (D))) */ ;
    defparam n30987_bdd_4_lut_4_lut_then_4_lut.init = 16'ha280;
    FD1P3AX block_reg_3___i1 (.D(write_data_c_0), .SP(clk_c_enable_2444), 
            .CK(clk_c), .Q(\block_reg[3] [0]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i1.GSR = "ENABLED";
    ROM256X1A sword_31__I_0_Mux_3 (.AD0(tmp_sboxw[24]), .AD1(tmp_sboxw[25]), 
            .AD2(tmp_sboxw[26]), .AD3(tmp_sboxw[27]), .AD4(tmp_sboxw[28]), 
            .AD5(tmp_sboxw[29]), .AD6(tmp_sboxw[30]), .AD7(tmp_sboxw[31]), 
            .DO0(new_sboxw_adj_9440[27])) /* synthesis initstate=0xC21A4F3CEDDCC8177B4DF9B4DA220CD1C67E14B661F51C623A33AB82E2758986 */ ;
    defparam sword_31__I_0_Mux_3.initval = 256'hC21A4F3CEDDCC8177B4DF9B4DA220CD1C67E14B661F51C623A33AB82E2758986;
    PFUMX i29066 (.BLUT(n34025), .ALUT(n34026), .C0(address_c_0), .Z(n34027));
    LUT4 n30987_bdd_4_lut_4_lut_else_4_lut (.A(n8904), .B(result_reg[87]), 
         .C(result_reg[119]), .D(address_c_0), .Z(n33962)) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam n30987_bdd_4_lut_4_lut_else_4_lut.init = 16'h88a0;
    PFUMX i29064 (.BLUT(n34022), .ALUT(n34023), .C0(address_c_0), .Z(n34024));
    ROM256X1A sword_31__I_0_Mux_5 (.AD0(tmp_sboxw[24]), .AD1(tmp_sboxw[25]), 
            .AD2(tmp_sboxw[26]), .AD3(tmp_sboxw[27]), .AD4(tmp_sboxw[28]), 
            .AD5(tmp_sboxw[29]), .AD6(tmp_sboxw[30]), .AD7(tmp_sboxw[31]), 
            .DO0(new_sboxw_adj_9440[29])) /* synthesis initstate=0xABBA8EF7872D518C98C5572AAF7EF2A1862233241073622F95DE21DA4167A5F4 */ ;
    defparam sword_31__I_0_Mux_5.initval = 256'hABBA8EF7872D518C98C5572AAF7EF2A1862233241073622F95DE21DA4167A5F4;
    ROM256X1A sword_31__I_0_Mux_6 (.AD0(tmp_sboxw[24]), .AD1(tmp_sboxw[25]), 
            .AD2(tmp_sboxw[26]), .AD3(tmp_sboxw[27]), .AD4(tmp_sboxw[28]), 
            .AD5(tmp_sboxw[29]), .AD6(tmp_sboxw[30]), .AD7(tmp_sboxw[31]), 
            .DO0(new_sboxw_adj_9440[30])) /* synthesis initstate=0x9B68A34AA647C842FE7B054BEB14DEF8811147420DBF3D2F5B28F323FC43E20D */ ;
    defparam sword_31__I_0_Mux_6.initval = 256'h9B68A34AA647C842FE7B054BEB14DEF8811147420DBF3D2F5B28F323FC43E20D;
    ROM256X1A sword_31__I_0_Mux_7 (.AD0(tmp_sboxw[24]), .AD1(tmp_sboxw[25]), 
            .AD2(tmp_sboxw[26]), .AD3(tmp_sboxw[27]), .AD4(tmp_sboxw[28]), 
            .AD5(tmp_sboxw[29]), .AD6(tmp_sboxw[30]), .AD7(tmp_sboxw[31]), 
            .DO0(new_sboxw_adj_9440[31])) /* synthesis initstate=0x015057D3FA286156AF3152C24BB37FC247193377F0F0CB5664A46534F2DAFD48 */ ;
    defparam sword_31__I_0_Mux_7.initval = 256'h015057D3FA286156AF3152C24BB37FC247193377F0F0CB5664A46534F2DAFD48;
    ROM256X1A sword_23__I_0_Mux_1 (.AD0(tmp_sboxw[16]), .AD1(tmp_sboxw[17]), 
            .AD2(tmp_sboxw[18]), .AD3(tmp_sboxw[19]), .AD4(tmp_sboxw[20]), 
            .AD5(tmp_sboxw[21]), .AD6(tmp_sboxw[22]), .AD7(tmp_sboxw[23]), 
            .DO0(new_sboxw_adj_9440[17])) /* synthesis initstate=0x08FB36349C4492694B3EDF05C519CFB1EAFCA1C41D80C095278AF97AA6FAED25 */ ;
    defparam sword_23__I_0_Mux_1.initval = 256'h08FB36349C4492694B3EDF05C519CFB1EAFCA1C41D80C095278AF97AA6FAED25;
    ROM256X1A sword_23__I_0_Mux_2 (.AD0(tmp_sboxw[16]), .AD1(tmp_sboxw[17]), 
            .AD2(tmp_sboxw[18]), .AD3(tmp_sboxw[19]), .AD4(tmp_sboxw[20]), 
            .AD5(tmp_sboxw[21]), .AD6(tmp_sboxw[22]), .AD7(tmp_sboxw[23]), 
            .DO0(new_sboxw_adj_9440[18])) /* synthesis initstate=0xD4ED0858CBA4D063A8174B51F4F76D70066ECB30FF317F9C914A87953BE14968 */ ;
    defparam sword_23__I_0_Mux_2.initval = 256'hD4ED0858CBA4D063A8174B51F4F76D70066ECB30FF317F9C914A87953BE14968;
    ROM256X1A sword_23__I_0_Mux_3 (.AD0(tmp_sboxw[16]), .AD1(tmp_sboxw[17]), 
            .AD2(tmp_sboxw[18]), .AD3(tmp_sboxw[19]), .AD4(tmp_sboxw[20]), 
            .AD5(tmp_sboxw[21]), .AD6(tmp_sboxw[22]), .AD7(tmp_sboxw[23]), 
            .DO0(new_sboxw_adj_9440[19])) /* synthesis initstate=0xC21A4F3CEDDCC8177B4DF9B4DA220CD1C67E14B661F51C623A33AB82E2758986 */ ;
    defparam sword_23__I_0_Mux_3.initval = 256'hC21A4F3CEDDCC8177B4DF9B4DA220CD1C67E14B661F51C623A33AB82E2758986;
    ROM256X1A sword_23__I_0_Mux_4 (.AD0(tmp_sboxw[16]), .AD1(tmp_sboxw[17]), 
            .AD2(tmp_sboxw[18]), .AD3(tmp_sboxw[19]), .AD4(tmp_sboxw[20]), 
            .AD5(tmp_sboxw[21]), .AD6(tmp_sboxw[22]), .AD7(tmp_sboxw[23]), 
            .DO0(new_sboxw_adj_9440[20])) /* synthesis initstate=0x94796CC45C368F8BDB67E21E7645B347242535634BDAD5C743A0248F2155E9B9 */ ;
    defparam sword_23__I_0_Mux_4.initval = 256'h94796CC45C368F8BDB67E21E7645B347242535634BDAD5C743A0248F2155E9B9;
    ROM256X1A sword_23__I_0_Mux_5 (.AD0(tmp_sboxw[16]), .AD1(tmp_sboxw[17]), 
            .AD2(tmp_sboxw[18]), .AD3(tmp_sboxw[19]), .AD4(tmp_sboxw[20]), 
            .AD5(tmp_sboxw[21]), .AD6(tmp_sboxw[22]), .AD7(tmp_sboxw[23]), 
            .DO0(new_sboxw_adj_9440[21])) /* synthesis initstate=0xABBA8EF7872D518C98C5572AAF7EF2A1862233241073622F95DE21DA4167A5F4 */ ;
    defparam sword_23__I_0_Mux_5.initval = 256'hABBA8EF7872D518C98C5572AAF7EF2A1862233241073622F95DE21DA4167A5F4;
    ROM256X1A sword_23__I_0_Mux_6 (.AD0(tmp_sboxw[16]), .AD1(tmp_sboxw[17]), 
            .AD2(tmp_sboxw[18]), .AD3(tmp_sboxw[19]), .AD4(tmp_sboxw[20]), 
            .AD5(tmp_sboxw[21]), .AD6(tmp_sboxw[22]), .AD7(tmp_sboxw[23]), 
            .DO0(new_sboxw_adj_9440[22])) /* synthesis initstate=0x9B68A34AA647C842FE7B054BEB14DEF8811147420DBF3D2F5B28F323FC43E20D */ ;
    defparam sword_23__I_0_Mux_6.initval = 256'h9B68A34AA647C842FE7B054BEB14DEF8811147420DBF3D2F5B28F323FC43E20D;
    ROM256X1A sword_23__I_0_Mux_7 (.AD0(tmp_sboxw[16]), .AD1(tmp_sboxw[17]), 
            .AD2(tmp_sboxw[18]), .AD3(tmp_sboxw[19]), .AD4(tmp_sboxw[20]), 
            .AD5(tmp_sboxw[21]), .AD6(tmp_sboxw[22]), .AD7(tmp_sboxw[23]), 
            .DO0(new_sboxw_adj_9440[23])) /* synthesis initstate=0x015057D3FA286156AF3152C24BB37FC247193377F0F0CB5664A46534F2DAFD48 */ ;
    defparam sword_23__I_0_Mux_7.initval = 256'h015057D3FA286156AF3152C24BB37FC247193377F0F0CB5664A46534F2DAFD48;
    ROM256X1A sword_15__I_0_Mux_1 (.AD0(tmp_sboxw[8]), .AD1(tmp_sboxw[9]), 
            .AD2(tmp_sboxw[10]), .AD3(tmp_sboxw[11]), .AD4(tmp_sboxw[12]), 
            .AD5(tmp_sboxw[13]), .AD6(tmp_sboxw[14]), .AD7(tmp_sboxw[15]), 
            .DO0(new_sboxw_adj_9440[9])) /* synthesis initstate=0x08FB36349C4492694B3EDF05C519CFB1EAFCA1C41D80C095278AF97AA6FAED25 */ ;
    defparam sword_15__I_0_Mux_1.initval = 256'h08FB36349C4492694B3EDF05C519CFB1EAFCA1C41D80C095278AF97AA6FAED25;
    ROM256X1A sword_15__I_0_Mux_2 (.AD0(tmp_sboxw[8]), .AD1(tmp_sboxw[9]), 
            .AD2(tmp_sboxw[10]), .AD3(tmp_sboxw[11]), .AD4(tmp_sboxw[12]), 
            .AD5(tmp_sboxw[13]), .AD6(tmp_sboxw[14]), .AD7(tmp_sboxw[15]), 
            .DO0(new_sboxw_adj_9440[10])) /* synthesis initstate=0xD4ED0858CBA4D063A8174B51F4F76D70066ECB30FF317F9C914A87953BE14968 */ ;
    defparam sword_15__I_0_Mux_2.initval = 256'hD4ED0858CBA4D063A8174B51F4F76D70066ECB30FF317F9C914A87953BE14968;
    ROM256X1A sword_15__I_0_Mux_3 (.AD0(tmp_sboxw[8]), .AD1(tmp_sboxw[9]), 
            .AD2(tmp_sboxw[10]), .AD3(tmp_sboxw[11]), .AD4(tmp_sboxw[12]), 
            .AD5(tmp_sboxw[13]), .AD6(tmp_sboxw[14]), .AD7(tmp_sboxw[15]), 
            .DO0(new_sboxw_adj_9440[11])) /* synthesis initstate=0xC21A4F3CEDDCC8177B4DF9B4DA220CD1C67E14B661F51C623A33AB82E2758986 */ ;
    defparam sword_15__I_0_Mux_3.initval = 256'hC21A4F3CEDDCC8177B4DF9B4DA220CD1C67E14B661F51C623A33AB82E2758986;
    ROM256X1A sword_15__I_0_Mux_4 (.AD0(tmp_sboxw[8]), .AD1(tmp_sboxw[9]), 
            .AD2(tmp_sboxw[10]), .AD3(tmp_sboxw[11]), .AD4(tmp_sboxw[12]), 
            .AD5(tmp_sboxw[13]), .AD6(tmp_sboxw[14]), .AD7(tmp_sboxw[15]), 
            .DO0(new_sboxw_adj_9440[12])) /* synthesis initstate=0x94796CC45C368F8BDB67E21E7645B347242535634BDAD5C743A0248F2155E9B9 */ ;
    defparam sword_15__I_0_Mux_4.initval = 256'h94796CC45C368F8BDB67E21E7645B347242535634BDAD5C743A0248F2155E9B9;
    ROM256X1A sword_15__I_0_Mux_5 (.AD0(tmp_sboxw[8]), .AD1(tmp_sboxw[9]), 
            .AD2(tmp_sboxw[10]), .AD3(tmp_sboxw[11]), .AD4(tmp_sboxw[12]), 
            .AD5(tmp_sboxw[13]), .AD6(tmp_sboxw[14]), .AD7(tmp_sboxw[15]), 
            .DO0(new_sboxw_adj_9440[13])) /* synthesis initstate=0xABBA8EF7872D518C98C5572AAF7EF2A1862233241073622F95DE21DA4167A5F4 */ ;
    defparam sword_15__I_0_Mux_5.initval = 256'hABBA8EF7872D518C98C5572AAF7EF2A1862233241073622F95DE21DA4167A5F4;
    ROM256X1A sword_15__I_0_Mux_6 (.AD0(tmp_sboxw[8]), .AD1(tmp_sboxw[9]), 
            .AD2(tmp_sboxw[10]), .AD3(tmp_sboxw[11]), .AD4(tmp_sboxw[12]), 
            .AD5(tmp_sboxw[13]), .AD6(tmp_sboxw[14]), .AD7(tmp_sboxw[15]), 
            .DO0(new_sboxw_adj_9440[14])) /* synthesis initstate=0x9B68A34AA647C842FE7B054BEB14DEF8811147420DBF3D2F5B28F323FC43E20D */ ;
    defparam sword_15__I_0_Mux_6.initval = 256'h9B68A34AA647C842FE7B054BEB14DEF8811147420DBF3D2F5B28F323FC43E20D;
    ROM256X1A sword_15__I_0_Mux_7 (.AD0(tmp_sboxw[8]), .AD1(tmp_sboxw[9]), 
            .AD2(tmp_sboxw[10]), .AD3(tmp_sboxw[11]), .AD4(tmp_sboxw[12]), 
            .AD5(tmp_sboxw[13]), .AD6(tmp_sboxw[14]), .AD7(tmp_sboxw[15]), 
            .DO0(new_sboxw_adj_9440[15])) /* synthesis initstate=0x015057D3FA286156AF3152C24BB37FC247193377F0F0CB5664A46534F2DAFD48 */ ;
    defparam sword_15__I_0_Mux_7.initval = 256'h015057D3FA286156AF3152C24BB37FC247193377F0F0CB5664A46534F2DAFD48;
    ROM256X1A sword_7__I_0_Mux_1 (.AD0(tmp_sboxw[0]), .AD1(tmp_sboxw[1]), 
            .AD2(tmp_sboxw[2]), .AD3(tmp_sboxw[3]), .AD4(tmp_sboxw[4]), 
            .AD5(tmp_sboxw[5]), .AD6(tmp_sboxw[6]), .AD7(tmp_sboxw[7]), 
            .DO0(new_sboxw_adj_9440[1])) /* synthesis initstate=0x08FB36349C4492694B3EDF05C519CFB1EAFCA1C41D80C095278AF97AA6FAED25 */ ;
    defparam sword_7__I_0_Mux_1.initval = 256'h08FB36349C4492694B3EDF05C519CFB1EAFCA1C41D80C095278AF97AA6FAED25;
    ROM256X1A sword_7__I_0_Mux_2 (.AD0(tmp_sboxw[0]), .AD1(tmp_sboxw[1]), 
            .AD2(tmp_sboxw[2]), .AD3(tmp_sboxw[3]), .AD4(tmp_sboxw[4]), 
            .AD5(tmp_sboxw[5]), .AD6(tmp_sboxw[6]), .AD7(tmp_sboxw[7]), 
            .DO0(new_sboxw_adj_9440[2])) /* synthesis initstate=0xD4ED0858CBA4D063A8174B51F4F76D70066ECB30FF317F9C914A87953BE14968 */ ;
    defparam sword_7__I_0_Mux_2.initval = 256'hD4ED0858CBA4D063A8174B51F4F76D70066ECB30FF317F9C914A87953BE14968;
    ROM256X1A sword_7__I_0_Mux_3 (.AD0(tmp_sboxw[0]), .AD1(tmp_sboxw[1]), 
            .AD2(tmp_sboxw[2]), .AD3(tmp_sboxw[3]), .AD4(tmp_sboxw[4]), 
            .AD5(tmp_sboxw[5]), .AD6(tmp_sboxw[6]), .AD7(tmp_sboxw[7]), 
            .DO0(new_sboxw_adj_9440[3])) /* synthesis initstate=0xC21A4F3CEDDCC8177B4DF9B4DA220CD1C67E14B661F51C623A33AB82E2758986 */ ;
    defparam sword_7__I_0_Mux_3.initval = 256'hC21A4F3CEDDCC8177B4DF9B4DA220CD1C67E14B661F51C623A33AB82E2758986;
    ROM256X1A sword_7__I_0_Mux_4 (.AD0(tmp_sboxw[0]), .AD1(tmp_sboxw[1]), 
            .AD2(tmp_sboxw[2]), .AD3(tmp_sboxw[3]), .AD4(tmp_sboxw[4]), 
            .AD5(tmp_sboxw[5]), .AD6(tmp_sboxw[6]), .AD7(tmp_sboxw[7]), 
            .DO0(new_sboxw_adj_9440[4])) /* synthesis initstate=0x94796CC45C368F8BDB67E21E7645B347242535634BDAD5C743A0248F2155E9B9 */ ;
    defparam sword_7__I_0_Mux_4.initval = 256'h94796CC45C368F8BDB67E21E7645B347242535634BDAD5C743A0248F2155E9B9;
    ROM256X1A sword_7__I_0_Mux_5 (.AD0(tmp_sboxw[0]), .AD1(tmp_sboxw[1]), 
            .AD2(tmp_sboxw[2]), .AD3(tmp_sboxw[3]), .AD4(tmp_sboxw[4]), 
            .AD5(tmp_sboxw[5]), .AD6(tmp_sboxw[6]), .AD7(tmp_sboxw[7]), 
            .DO0(new_sboxw_adj_9440[5])) /* synthesis initstate=0xABBA8EF7872D518C98C5572AAF7EF2A1862233241073622F95DE21DA4167A5F4 */ ;
    defparam sword_7__I_0_Mux_5.initval = 256'hABBA8EF7872D518C98C5572AAF7EF2A1862233241073622F95DE21DA4167A5F4;
    ROM256X1A sword_7__I_0_Mux_6 (.AD0(tmp_sboxw[0]), .AD1(tmp_sboxw[1]), 
            .AD2(tmp_sboxw[2]), .AD3(tmp_sboxw[3]), .AD4(tmp_sboxw[4]), 
            .AD5(tmp_sboxw[5]), .AD6(tmp_sboxw[6]), .AD7(tmp_sboxw[7]), 
            .DO0(new_sboxw_adj_9440[6])) /* synthesis initstate=0x9B68A34AA647C842FE7B054BEB14DEF8811147420DBF3D2F5B28F323FC43E20D */ ;
    defparam sword_7__I_0_Mux_6.initval = 256'h9B68A34AA647C842FE7B054BEB14DEF8811147420DBF3D2F5B28F323FC43E20D;
    ROM256X1A sword_7__I_0_Mux_7 (.AD0(tmp_sboxw[0]), .AD1(tmp_sboxw[1]), 
            .AD2(tmp_sboxw[2]), .AD3(tmp_sboxw[3]), .AD4(tmp_sboxw[4]), 
            .AD5(tmp_sboxw[5]), .AD6(tmp_sboxw[6]), .AD7(tmp_sboxw[7]), 
            .DO0(new_sboxw_adj_9440[7])) /* synthesis initstate=0x015057D3FA286156AF3152C24BB37FC247193377F0F0CB5664A46534F2DAFD48 */ ;
    defparam sword_7__I_0_Mux_7.initval = 256'h015057D3FA286156AF3152C24BB37FC247193377F0F0CB5664A46534F2DAFD48;
    ROM256X1A sword_7__I_0_Mux_0 (.AD0(tmp_sboxw[0]), .AD1(tmp_sboxw[1]), 
            .AD2(tmp_sboxw[2]), .AD3(tmp_sboxw[3]), .AD4(tmp_sboxw[4]), 
            .AD5(tmp_sboxw[5]), .AD6(tmp_sboxw[6]), .AD7(tmp_sboxw[7]), 
            .DO0(new_sboxw_adj_9440[0])) /* synthesis initstate=0xBB23F64CBBBE99EB224883FB66F0853EBF6869447A703000FA244CC2C4F6F54A */ ;
    defparam sword_7__I_0_Mux_0.initval = 256'hBB23F64CBBBE99EB224883FB66F0853EBF6869447A703000FA244CC2C4F6F54A;
    ROM256X1A sword_15__I_0_Mux_0 (.AD0(tmp_sboxw[8]), .AD1(tmp_sboxw[9]), 
            .AD2(tmp_sboxw[10]), .AD3(tmp_sboxw[11]), .AD4(tmp_sboxw[12]), 
            .AD5(tmp_sboxw[13]), .AD6(tmp_sboxw[14]), .AD7(tmp_sboxw[15]), 
            .DO0(new_sboxw_adj_9440[8])) /* synthesis initstate=0xBB23F64CBBBE99EB224883FB66F0853EBF6869447A703000FA244CC2C4F6F54A */ ;
    defparam sword_15__I_0_Mux_0.initval = 256'hBB23F64CBBBE99EB224883FB66F0853EBF6869447A703000FA244CC2C4F6F54A;
    ROM256X1A sword_23__I_0_Mux_0 (.AD0(tmp_sboxw[16]), .AD1(tmp_sboxw[17]), 
            .AD2(tmp_sboxw[18]), .AD3(tmp_sboxw[19]), .AD4(tmp_sboxw[20]), 
            .AD5(tmp_sboxw[21]), .AD6(tmp_sboxw[22]), .AD7(tmp_sboxw[23]), 
            .DO0(new_sboxw_adj_9440[16])) /* synthesis initstate=0xBB23F64CBBBE99EB224883FB66F0853EBF6869447A703000FA244CC2C4F6F54A */ ;
    defparam sword_23__I_0_Mux_0.initval = 256'hBB23F64CBBBE99EB224883FB66F0853EBF6869447A703000FA244CC2C4F6F54A;
    ROM256X1A sword_31__I_0_Mux_0 (.AD0(tmp_sboxw[24]), .AD1(tmp_sboxw[25]), 
            .AD2(tmp_sboxw[26]), .AD3(tmp_sboxw[27]), .AD4(tmp_sboxw[28]), 
            .AD5(tmp_sboxw[29]), .AD6(tmp_sboxw[30]), .AD7(tmp_sboxw[31]), 
            .DO0(new_sboxw_adj_9440[24])) /* synthesis initstate=0xBB23F64CBBBE99EB224883FB66F0853EBF6869447A703000FA244CC2C4F6F54A */ ;
    defparam sword_31__I_0_Mux_0.initval = 256'hBB23F64CBBBE99EB224883FB66F0853EBF6869447A703000FA244CC2C4F6F54A;
    ROM256X1A sboxw_23__I_0_Mux_0 (.AD0(muxed_sboxw[16]), .AD1(muxed_sboxw[17]), 
            .AD2(muxed_sboxw[18]), .AD3(muxed_sboxw[19]), .AD4(muxed_sboxw[20]), 
            .AD5(muxed_sboxw[21]), .AD6(muxed_sboxw[22]), .AD7(muxed_sboxw[23]), 
            .DO0(new_sboxw[16])) /* synthesis initstate=0x4F1EAD396F247A0410BDB210C006EAB568AB4BFA8ACB7A13B14EDE67096C6EED */ ;
    defparam sboxw_23__I_0_Mux_0.initval = 256'h4F1EAD396F247A0410BDB210C006EAB568AB4BFA8ACB7A13B14EDE67096C6EED;
    ROM256X1A sboxw_23__I_0_Mux_1 (.AD0(muxed_sboxw[16]), .AD1(muxed_sboxw[17]), 
            .AD2(muxed_sboxw[18]), .AD3(muxed_sboxw[19]), .AD4(muxed_sboxw[20]), 
            .AD5(muxed_sboxw[21]), .AD6(muxed_sboxw[22]), .AD7(muxed_sboxw[23]), 
            .DO0(new_sboxw[17])) /* synthesis initstate=0xC870974094EAD8A96A450B2EF33486B4E61A4C5E97816F7A7BAE007D4C53FC7D */ ;
    defparam sboxw_23__I_0_Mux_1.initval = 256'hC870974094EAD8A96A450B2EF33486B4E61A4C5E97816F7A7BAE007D4C53FC7D;
    ROM256X1A sboxw_23__I_0_Mux_2 (.AD0(muxed_sboxw[16]), .AD1(muxed_sboxw[17]), 
            .AD2(muxed_sboxw[18]), .AD3(muxed_sboxw[19]), .AD4(muxed_sboxw[20]), 
            .AD5(muxed_sboxw[21]), .AD6(muxed_sboxw[22]), .AD7(muxed_sboxw[23]), 
            .DO0(new_sboxw[18])) /* synthesis initstate=0xAC39B6C0D6CE2EFC577D64E03B0C3FFB23A869A2A428C424A16387FB3B48B4C6 */ ;
    defparam sboxw_23__I_0_Mux_2.initval = 256'hAC39B6C0D6CE2EFC577D64E03B0C3FFB23A869A2A428C424A16387FB3B48B4C6;
    ROM256X1A sboxw_23__I_0_Mux_3 (.AD0(muxed_sboxw[16]), .AD1(muxed_sboxw[17]), 
            .AD2(muxed_sboxw[18]), .AD3(muxed_sboxw[19]), .AD4(muxed_sboxw[20]), 
            .AD5(muxed_sboxw[21]), .AD6(muxed_sboxw[22]), .AD7(muxed_sboxw[23]), 
            .DO0(new_sboxw[19])) /* synthesis initstate=0x4E9DDB76C892FB1BE9DA849CF6AC6C1B2568EA2EFFA8527D109020A2193D586A */ ;
    defparam sboxw_23__I_0_Mux_3.initval = 256'h4E9DDB76C892FB1BE9DA849CF6AC6C1B2568EA2EFFA8527D109020A2193D586A;
    ROM256X1A sboxw_23__I_0_Mux_4 (.AD0(muxed_sboxw[16]), .AD1(muxed_sboxw[17]), 
            .AD2(muxed_sboxw[18]), .AD3(muxed_sboxw[19]), .AD4(muxed_sboxw[20]), 
            .AD5(muxed_sboxw[21]), .AD6(muxed_sboxw[22]), .AD7(muxed_sboxw[23]), 
            .DO0(new_sboxw[20])) /* synthesis initstate=0xF210A3AECE472E532624B286BC48ECB4F7F17A494CE30F58C2B0F97752B8B11E */ ;
    defparam sboxw_23__I_0_Mux_4.initval = 256'hF210A3AECE472E532624B286BC48ECB4F7F17A494CE30F58C2B0F97752B8B11E;
    ROM256X1A sboxw_23__I_0_Mux_5 (.AD0(muxed_sboxw[16]), .AD1(muxed_sboxw[17]), 
            .AD2(muxed_sboxw[18]), .AD3(muxed_sboxw[19]), .AD4(muxed_sboxw[20]), 
            .AD5(muxed_sboxw[21]), .AD6(muxed_sboxw[22]), .AD7(muxed_sboxw[23]), 
            .DO0(new_sboxw[21])) /* synthesis initstate=0x54B248130B4F256F7D8DCC4706319E086BC2AA4E0D787AA4F8045F7B6D98DD7F */ ;
    defparam sboxw_23__I_0_Mux_5.initval = 256'h54B248130B4F256F7D8DCC4706319E086BC2AA4E0D787AA4F8045F7B6D98DD7F;
    ROM256X1A sboxw_23__I_0_Mux_6 (.AD0(muxed_sboxw[16]), .AD1(muxed_sboxw[17]), 
            .AD2(muxed_sboxw[18]), .AD3(muxed_sboxw[19]), .AD4(muxed_sboxw[20]), 
            .AD5(muxed_sboxw[21]), .AD6(muxed_sboxw[22]), .AD7(muxed_sboxw[23]), 
            .DO0(new_sboxw[22])) /* synthesis initstate=0x21E0B833255917823F6BCB91B30DB559E4851B3BF3AB2560980A3CC2C2FDB4FF */ ;
    defparam sboxw_23__I_0_Mux_6.initval = 256'h21E0B833255917823F6BCB91B30DB559E4851B3BF3AB2560980A3CC2C2FDB4FF;
    ROM256X1A sword_31__I_0_Mux_4 (.AD0(tmp_sboxw[24]), .AD1(tmp_sboxw[25]), 
            .AD2(tmp_sboxw[26]), .AD3(tmp_sboxw[27]), .AD4(tmp_sboxw[28]), 
            .AD5(tmp_sboxw[29]), .AD6(tmp_sboxw[30]), .AD7(tmp_sboxw[31]), 
            .DO0(new_sboxw_adj_9440[28])) /* synthesis initstate=0x94796CC45C368F8BDB67E21E7645B347242535634BDAD5C743A0248F2155E9B9 */ ;
    defparam sword_31__I_0_Mux_4.initval = 256'h94796CC45C368F8BDB67E21E7645B347242535634BDAD5C743A0248F2155E9B9;
    ROM256X1A sboxw_23__I_0_Mux_7 (.AD0(muxed_sboxw[16]), .AD1(muxed_sboxw[17]), 
            .AD2(muxed_sboxw[18]), .AD3(muxed_sboxw[19]), .AD4(muxed_sboxw[20]), 
            .AD5(muxed_sboxw[21]), .AD6(muxed_sboxw[22]), .AD7(muxed_sboxw[23]), 
            .DO0(new_sboxw[23])) /* synthesis initstate=0x52379DE7B844E3E14CB3770196CA0329E7BAC28F866AAC825CAA2EC7BF977090 */ ;
    defparam sboxw_23__I_0_Mux_7.initval = 256'h52379DE7B844E3E14CB3770196CA0329E7BAC28F866AAC825CAA2EC7BF977090;
    ROM256X1A sword_31__I_0_Mux_1 (.AD0(tmp_sboxw[24]), .AD1(tmp_sboxw[25]), 
            .AD2(tmp_sboxw[26]), .AD3(tmp_sboxw[27]), .AD4(tmp_sboxw[28]), 
            .AD5(tmp_sboxw[29]), .AD6(tmp_sboxw[30]), .AD7(tmp_sboxw[31]), 
            .DO0(new_sboxw_adj_9440[25])) /* synthesis initstate=0x08FB36349C4492694B3EDF05C519CFB1EAFCA1C41D80C095278AF97AA6FAED25 */ ;
    defparam sword_31__I_0_Mux_1.initval = 256'h08FB36349C4492694B3EDF05C519CFB1EAFCA1C41D80C095278AF97AA6FAED25;
    ROM256X1A sword_31__I_0_Mux_2 (.AD0(tmp_sboxw[24]), .AD1(tmp_sboxw[25]), 
            .AD2(tmp_sboxw[26]), .AD3(tmp_sboxw[27]), .AD4(tmp_sboxw[28]), 
            .AD5(tmp_sboxw[29]), .AD6(tmp_sboxw[30]), .AD7(tmp_sboxw[31]), 
            .DO0(new_sboxw_adj_9440[26])) /* synthesis initstate=0xD4ED0858CBA4D063A8174B51F4F76D70066ECB30FF317F9C914A87953BE14968 */ ;
    defparam sword_31__I_0_Mux_2.initval = 256'hD4ED0858CBA4D063A8174B51F4F76D70066ECB30FF317F9C914A87953BE14968;
    LUT4 i14937_4_lut (.A(n37), .B(n33950), .C(n34042), .D(n1504), .Z(read_data_c_30)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B+!(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(249[13] 264[16])
    defparam i14937_4_lut.init = 16'h3011;
    LUT4 i2_4_lut (.A(address_c_3), .B(address_c_4), .C(address_c_2), 
         .D(n28824), .Z(n1504)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i2_4_lut.init = 16'h0400;
    PFUMX i29062 (.BLUT(n34019), .ALUT(n34020), .C0(address_c_0), .Z(n34021));
    OB read_data_pad_30 (.I(read_data_c_30), .O(read_data[30]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(51[33:42])
    OB read_data_pad_31 (.I(read_data_c_31), .O(read_data[31]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(51[33:42])
    LUT4 n30978_bdd_4_lut_4_lut_then_4_lut (.A(n8904), .B(address_c_0), 
         .C(result_reg[20]), .D(result_reg[52]), .Z(n33954)) /* synthesis lut_function=(A (B (C)+!B (D))) */ ;
    defparam n30978_bdd_4_lut_4_lut_then_4_lut.init = 16'ha280;
    LUT4 n30978_bdd_4_lut_4_lut_else_4_lut (.A(n8904), .B(result_reg[84]), 
         .C(result_reg[116]), .D(address_c_0), .Z(n33953)) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam n30978_bdd_4_lut_4_lut_else_4_lut.init = 16'h88a0;
    FD1P3AX encdec_reg_105 (.D(write_data_c_0), .SP(config_we), .CK(clk_c), 
            .Q(encdec_reg));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam encdec_reg_105.GSR = "ENABLED";
    FD1P3AX keylen_reg_106 (.D(write_data_c_1), .SP(config_we), .CK(clk_c), 
            .Q(\key_mem_ctrl.num_rounds [2]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam keylen_reg_106.GSR = "ENABLED";
    LUT4 i14936_4_lut (.A(n25954), .B(n33950), .C(n34039), .D(n1504), 
         .Z(read_data_c_29)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B+!(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(249[13] 264[16])
    defparam i14936_4_lut.init = 16'h3011;
    LUT4 i14935_4_lut (.A(n33), .B(n33950), .C(n34036), .D(n1504), .Z(read_data_c_28)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B+!(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(249[13] 264[16])
    defparam i14935_4_lut.init = 16'h3011;
    LUT4 i14934_4_lut (.A(n37), .B(n33950), .C(n34033), .D(n1504), .Z(read_data_c_24)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B+!(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(249[13] 264[16])
    defparam i14934_4_lut.init = 16'h3011;
    PFUMX i29060 (.BLUT(n34016), .ALUT(n34017), .C0(address_c_0), .Z(n34018));
    LUT4 i14933_4_lut (.A(n37), .B(n33950), .C(n34030), .D(n1504), .Z(read_data_c_22)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B+!(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(249[13] 264[16])
    defparam i14933_4_lut.init = 16'h3011;
    LUT4 i14932_4_lut (.A(n25954), .B(n33950), .C(n34027), .D(n1504), 
         .Z(read_data_c_21)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B+!(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(249[13] 264[16])
    defparam i14932_4_lut.init = 16'h3011;
    LUT4 i14931_4_lut (.A(n33), .B(n33950), .C(n34024), .D(n1504), .Z(read_data_c_19)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B+!(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(249[13] 264[16])
    defparam i14931_4_lut.init = 16'h3011;
    LUT4 i14930_4_lut (.A(n20756), .B(n33950), .C(n34021), .D(n1504), 
         .Z(read_data_c_18)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B+!(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(249[13] 264[16])
    defparam i14930_4_lut.init = 16'h3011;
    LUT4 i14929_4_lut (.A(n33), .B(n33950), .C(n34018), .D(n1504), .Z(read_data_c_17)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B+!(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(249[13] 264[16])
    defparam i14929_4_lut.init = 16'h3011;
    LUT4 i14928_4_lut (.A(n37), .B(n33950), .C(n34015), .D(n1504), .Z(read_data_c_16)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B+!(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(249[13] 264[16])
    defparam i14928_4_lut.init = 16'h3011;
    LUT4 i14927_4_lut (.A(n37), .B(n33950), .C(n34012), .D(n1504), .Z(read_data_c_14)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B+!(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(249[13] 264[16])
    defparam i14927_4_lut.init = 16'h3011;
    LUT4 i14926_4_lut (.A(n25954), .B(n33950), .C(n34009), .D(n1504), 
         .Z(read_data_c_13)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B+!(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(249[13] 264[16])
    defparam i14926_4_lut.init = 16'h3011;
    LUT4 i14925_4_lut (.A(n20756), .B(n33950), .C(n34006), .D(n1504), 
         .Z(read_data_c_12)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B+!(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(249[13] 264[16])
    defparam i14925_4_lut.init = 16'h3011;
    LUT4 i14924_4_lut (.A(n33), .B(n33950), .C(n34003), .D(n1504), .Z(read_data_c_10)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B+!(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(249[13] 264[16])
    defparam i14924_4_lut.init = 16'h3011;
    LUT4 i14923_4_lut (.A(n20756), .B(n33950), .C(n34000), .D(n1504), 
         .Z(read_data_c_9)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B+!(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(249[13] 264[16])
    defparam i14923_4_lut.init = 16'h3011;
    LUT4 i14922_4_lut (.A(n37), .B(n33950), .C(n33997), .D(n1504), .Z(read_data_c_8)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B+!(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(249[13] 264[16])
    defparam i14922_4_lut.init = 16'h3011;
    LUT4 i14921_4_lut (.A(n25954), .B(n33950), .C(n33994), .D(n1504), 
         .Z(read_data_c_5)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B+!(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(249[13] 264[16])
    defparam i14921_4_lut.init = 16'h3011;
    LUT4 i14920_4_lut (.A(n33), .B(n33950), .C(n33991), .D(n1504), .Z(read_data_c_4)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B+!(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(249[13] 264[16])
    defparam i14920_4_lut.init = 16'h3011;
    LUT4 i1_4_lut (.A(n28845), .B(n28841), .C(n34048), .D(n1504), .Z(read_data_c_3)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut.init = 16'hc088;
    LUT4 i1_2_lut (.A(cs_c), .B(we_c), .Z(n28841)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut.init = 16'h2222;
    LUT4 i1_4_lut_adj_843 (.A(n28846), .B(n28841), .C(n34045), .D(n1504), 
         .Z(read_data_c_2)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_843.init = 16'hc088;
    LUT4 i1_4_lut_adj_844 (.A(n33950), .B(n28832), .C(n33988), .D(n1504), 
         .Z(read_data_c_1)) /* synthesis lut_function=(!(A+!(B (C+!(D))+!B (C (D))))) */ ;
    defparam i1_4_lut_adj_844.init = 16'h5044;
    LUT4 i1_4_lut_adj_845 (.A(n28830), .B(aes_core_ctrl_new_1__N_858[1]), 
         .C(valid_reg), .D(address_c_0), .Z(n28832)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_845.init = 16'ha088;
    LUT4 i1_4_lut_adj_846 (.A(n33950), .B(n28831), .C(n33985), .D(n1504), 
         .Z(read_data_c_0)) /* synthesis lut_function=(!(A+!(B (C+!(D))+!B (C (D))))) */ ;
    defparam i1_4_lut_adj_846.init = 16'h5044;
    LUT4 i1_4_lut_adj_847 (.A(n28830), .B(key_mem_ctrl_new_2__N_4928[0]), 
         .C(ready_reg), .D(address_c_0), .Z(n28831)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_847.init = 16'ha088;
    PFUMX i29058 (.BLUT(n34013), .ALUT(n34014), .C0(address_c_0), .Z(n34015));
    PFUMX i29056 (.BLUT(n34010), .ALUT(n34011), .C0(address_c_0), .Z(n34012));
    LUT4 n30996_bdd_4_lut_4_lut_then_4_lut (.A(n8904), .B(address_c_0), 
         .C(result_reg[26]), .D(result_reg[58]), .Z(n33966)) /* synthesis lut_function=(A (B (C)+!B (D))) */ ;
    defparam n30996_bdd_4_lut_4_lut_then_4_lut.init = 16'ha280;
    LUT4 n30996_bdd_4_lut_4_lut_else_4_lut (.A(n8904), .B(result_reg[90]), 
         .C(result_reg[122]), .D(address_c_0), .Z(n33965)) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam n30996_bdd_4_lut_4_lut_else_4_lut.init = 16'h88a0;
    PFUMX i29054 (.BLUT(n34007), .ALUT(n34008), .C0(address_c_0), .Z(n34009));
    LUT4 n30939_bdd_4_lut_4_lut_then_4_lut (.A(n8904), .B(address_c_0), 
         .C(result_reg[7]), .D(result_reg[39]), .Z(n33969)) /* synthesis lut_function=(A (B (C)+!B (D))) */ ;
    defparam n30939_bdd_4_lut_4_lut_then_4_lut.init = 16'ha280;
    LUT4 n30939_bdd_4_lut_4_lut_else_4_lut (.A(n8904), .B(result_reg[71]), 
         .C(result_reg[103]), .D(address_c_0), .Z(n33968)) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam n30939_bdd_4_lut_4_lut_else_4_lut.init = 16'h88a0;
    LUT4 n31011_bdd_4_lut_4_lut_then_4_lut (.A(n8904), .B(address_c_0), 
         .C(result_reg[31]), .D(result_reg[63]), .Z(n33972)) /* synthesis lut_function=(A (B (C)+!B (D))) */ ;
    defparam n31011_bdd_4_lut_4_lut_then_4_lut.init = 16'ha280;
    LUT4 n31011_bdd_4_lut_4_lut_else_4_lut (.A(n8904), .B(result_reg[95]), 
         .C(result_reg[127]), .D(address_c_0), .Z(n33971)) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam n31011_bdd_4_lut_4_lut_else_4_lut.init = 16'h88a0;
    PFUMX i29052 (.BLUT(n34004), .ALUT(n34005), .C0(address_c_0), .Z(n34006));
    LUT4 n30993_bdd_4_lut_4_lut_then_4_lut (.A(n8904), .B(address_c_0), 
         .C(result_reg[25]), .D(result_reg[57]), .Z(n33975)) /* synthesis lut_function=(A (B (C)+!B (D))) */ ;
    defparam n30993_bdd_4_lut_4_lut_then_4_lut.init = 16'ha280;
    LUT4 n30993_bdd_4_lut_4_lut_else_4_lut (.A(n8904), .B(result_reg[89]), 
         .C(result_reg[121]), .D(address_c_0), .Z(n33974)) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam n30993_bdd_4_lut_4_lut_else_4_lut.init = 16'h88a0;
    LUT4 n30963_bdd_4_lut_4_lut_then_4_lut (.A(n8904), .B(address_c_0), 
         .C(result_reg[15]), .D(result_reg[47]), .Z(n33978)) /* synthesis lut_function=(A (B (C)+!B (D))) */ ;
    defparam n30963_bdd_4_lut_4_lut_then_4_lut.init = 16'ha280;
    LUT4 n30963_bdd_4_lut_4_lut_else_4_lut (.A(n8904), .B(result_reg[79]), 
         .C(result_reg[111]), .D(address_c_0), .Z(n33977)) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam n30963_bdd_4_lut_4_lut_else_4_lut.init = 16'h88a0;
    LUT4 n30999_bdd_4_lut_4_lut_then_4_lut (.A(n8904), .B(address_c_0), 
         .C(result_reg[27]), .D(result_reg[59]), .Z(n33981)) /* synthesis lut_function=(A (B (C)+!B (D))) */ ;
    defparam n30999_bdd_4_lut_4_lut_then_4_lut.init = 16'ha280;
    LUT4 n30999_bdd_4_lut_4_lut_else_4_lut (.A(n8904), .B(result_reg[91]), 
         .C(result_reg[123]), .D(address_c_0), .Z(n33980)) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam n30999_bdd_4_lut_4_lut_else_4_lut.init = 16'h88a0;
    LUT4 i25767_then_3_lut (.A(result_reg[64]), .B(address_c_1), .C(result_reg[0]), 
         .Z(n33984)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i25767_then_3_lut.init = 16'he2e2;
    LUT4 i25767_else_3_lut (.A(result_reg[96]), .B(address_c_1), .C(result_reg[32]), 
         .Z(n33983)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i25767_else_3_lut.init = 16'he2e2;
    LUT4 i27858_2_lut_3_lut_4_lut (.A(address_c_2), .B(n33850), .C(address_c_1), 
         .D(address_c_0), .Z(clk_c_enable_387)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i27858_2_lut_3_lut_4_lut.init = 16'h0004;
    LUT4 i27890_2_lut_3_lut_4_lut (.A(address_c_2), .B(n33850), .C(address_c_1), 
         .D(address_c_0), .Z(clk_c_enable_323)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i27890_2_lut_3_lut_4_lut.init = 16'h0040;
    LUT4 i1_2_lut_4_lut (.A(address_c_2), .B(address_c_0), .C(n33850), 
         .D(address_c_1), .Z(clk_c_enable_195)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(49[33:40])
    defparam i1_2_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_4_lut_adj_848 (.A(address_c_2), .B(address_c_0), .C(n33850), 
         .D(address_c_1), .Z(clk_c_enable_259)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(49[33:40])
    defparam i1_2_lut_4_lut_adj_848.init = 16'h0020;
    LUT4 i15234_2_lut_4_lut (.A(n33910), .B(n28824), .C(n33857), .D(n33941), 
         .Z(clk_c_enable_2444)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i15234_2_lut_4_lut.init = 16'h4000;
    LUT4 i25770_then_3_lut (.A(result_reg[65]), .B(address_c_1), .C(result_reg[1]), 
         .Z(n33987)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i25770_then_3_lut.init = 16'he2e2;
    LUT4 i25770_else_3_lut (.A(result_reg[97]), .B(address_c_1), .C(result_reg[33]), 
         .Z(n33986)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i25770_else_3_lut.init = 16'he2e2;
    LUT4 i25773_then_3_lut (.A(result_reg[68]), .B(address_c_1), .C(result_reg[4]), 
         .Z(n33990)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i25773_then_3_lut.init = 16'he2e2;
    LUT4 i25773_else_3_lut (.A(result_reg[100]), .B(address_c_1), .C(result_reg[36]), 
         .Z(n33989)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i25773_else_3_lut.init = 16'he2e2;
    LUT4 i1_2_lut_4_lut_adj_849 (.A(address_c_3), .B(n33861), .C(n33949), 
         .D(\key_mem_ctrl.num_rounds [2]), .Z(n28845)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_2_lut_4_lut_adj_849.init = 16'h0200;
    LUT4 i1_2_lut_4_lut_adj_850 (.A(address_c_3), .B(n33861), .C(n33949), 
         .D(encdec_reg), .Z(n28846)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_2_lut_4_lut_adj_850.init = 16'h0200;
    LUT4 i2_3_lut_4_lut (.A(address_c_3), .B(n33861), .C(n33939), .D(n33946), 
         .Z(config_we)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(49[33:40])
    defparam i2_3_lut_4_lut.init = 16'h0020;
    LUT4 i25776_then_3_lut (.A(result_reg[69]), .B(address_c_1), .C(result_reg[5]), 
         .Z(n33993)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i25776_then_3_lut.init = 16'he2e2;
    LUT4 i25776_else_3_lut (.A(result_reg[101]), .B(address_c_1), .C(result_reg[37]), 
         .Z(n33992)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i25776_else_3_lut.init = 16'he2e2;
    OB read_data_pad_29 (.I(read_data_c_29), .O(read_data[29]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(51[33:42])
    FD1S3AX result_reg_i27 (.D(core_result[27]), .CK(clk_c), .Q(result_reg[27]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i27.GSR = "ENABLED";
    OB read_data_pad_28 (.I(read_data_c_28), .O(read_data[28]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(51[33:42])
    OB read_data_pad_27 (.I(read_data_c_27), .O(read_data[27]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(51[33:42])
    OB read_data_pad_26 (.I(read_data_c_26), .O(read_data[26]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(51[33:42])
    OB read_data_pad_25 (.I(read_data_c_25), .O(read_data[25]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(51[33:42])
    OB read_data_pad_24 (.I(read_data_c_24), .O(read_data[24]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(51[33:42])
    OB read_data_pad_23 (.I(read_data_c_23), .O(read_data[23]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(51[33:42])
    OB read_data_pad_22 (.I(read_data_c_22), .O(read_data[22]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(51[33:42])
    OB read_data_pad_21 (.I(read_data_c_21), .O(read_data[21]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(51[33:42])
    OB read_data_pad_20 (.I(read_data_c_20), .O(read_data[20]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(51[33:42])
    OB read_data_pad_19 (.I(read_data_c_19), .O(read_data[19]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(51[33:42])
    OB read_data_pad_18 (.I(read_data_c_18), .O(read_data[18]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(51[33:42])
    OB read_data_pad_17 (.I(read_data_c_17), .O(read_data[17]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(51[33:42])
    OB read_data_pad_16 (.I(read_data_c_16), .O(read_data[16]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(51[33:42])
    OB read_data_pad_15 (.I(read_data_c_15), .O(read_data[15]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(51[33:42])
    OB read_data_pad_14 (.I(read_data_c_14), .O(read_data[14]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(51[33:42])
    OB read_data_pad_13 (.I(read_data_c_13), .O(read_data[13]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(51[33:42])
    OB read_data_pad_12 (.I(read_data_c_12), .O(read_data[12]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(51[33:42])
    OB read_data_pad_11 (.I(read_data_c_11), .O(read_data[11]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(51[33:42])
    OB read_data_pad_10 (.I(read_data_c_10), .O(read_data[10]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(51[33:42])
    OB read_data_pad_9 (.I(read_data_c_9), .O(read_data[9]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(51[33:42])
    OB read_data_pad_8 (.I(read_data_c_8), .O(read_data[8]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(51[33:42])
    OB read_data_pad_7 (.I(read_data_c_7), .O(read_data[7]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(51[33:42])
    OB read_data_pad_6 (.I(read_data_c_6), .O(read_data[6]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(51[33:42])
    OB read_data_pad_5 (.I(read_data_c_5), .O(read_data[5]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(51[33:42])
    OB read_data_pad_4 (.I(read_data_c_4), .O(read_data[4]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(51[33:42])
    OB read_data_pad_3 (.I(read_data_c_3), .O(read_data[3]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(51[33:42])
    OB read_data_pad_2 (.I(read_data_c_2), .O(read_data[2]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(51[33:42])
    OB read_data_pad_1 (.I(read_data_c_1), .O(read_data[1]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(51[33:42])
    OB read_data_pad_0 (.I(read_data_c_0), .O(read_data[0]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(51[33:42])
    IB clk_pad (.I(clk), .O(clk_c));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(41[33:36])
    IB reset_n_pad (.I(reset_n), .O(reset_n_c));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(42[33:40])
    IB cs_pad (.I(cs), .O(cs_c));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(45[33:35])
    IB we_pad (.I(we), .O(we_c));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(46[33:35])
    IB address_pad_7 (.I(address[7]), .O(address_c_7));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(49[33:40])
    IB address_pad_6 (.I(address[6]), .O(address_c_6));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(49[33:40])
    IB address_pad_5 (.I(address[5]), .O(address_c_5));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(49[33:40])
    IB address_pad_4 (.I(address[4]), .O(address_c_4));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(49[33:40])
    IB address_pad_3 (.I(address[3]), .O(address_c_3));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(49[33:40])
    IB address_pad_2 (.I(address[2]), .O(address_c_2));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(49[33:40])
    IB address_pad_1 (.I(address[1]), .O(address_c_1));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(49[33:40])
    IB address_pad_0 (.I(address[0]), .O(address_c_0));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(49[33:40])
    IB write_data_pad_31 (.I(write_data[31]), .O(write_data_c_31));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(50[33:43])
    IB write_data_pad_30 (.I(write_data[30]), .O(write_data_c_30));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(50[33:43])
    IB write_data_pad_29 (.I(write_data[29]), .O(write_data_c_29));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(50[33:43])
    IB write_data_pad_28 (.I(write_data[28]), .O(write_data_c_28));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(50[33:43])
    IB write_data_pad_27 (.I(write_data[27]), .O(write_data_c_27));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(50[33:43])
    IB write_data_pad_26 (.I(write_data[26]), .O(write_data_c_26));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(50[33:43])
    IB write_data_pad_25 (.I(write_data[25]), .O(write_data_c_25));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(50[33:43])
    IB write_data_pad_24 (.I(write_data[24]), .O(write_data_c_24));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(50[33:43])
    IB write_data_pad_23 (.I(write_data[23]), .O(write_data_c_23));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(50[33:43])
    IB write_data_pad_22 (.I(write_data[22]), .O(write_data_c_22));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(50[33:43])
    IB write_data_pad_21 (.I(write_data[21]), .O(write_data_c_21));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(50[33:43])
    IB write_data_pad_20 (.I(write_data[20]), .O(write_data_c_20));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(50[33:43])
    IB write_data_pad_19 (.I(write_data[19]), .O(write_data_c_19));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(50[33:43])
    IB write_data_pad_18 (.I(write_data[18]), .O(write_data_c_18));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(50[33:43])
    IB write_data_pad_17 (.I(write_data[17]), .O(write_data_c_17));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(50[33:43])
    IB write_data_pad_16 (.I(write_data[16]), .O(write_data_c_16));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(50[33:43])
    IB write_data_pad_15 (.I(write_data[15]), .O(write_data_c_15));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(50[33:43])
    IB write_data_pad_14 (.I(write_data[14]), .O(write_data_c_14));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(50[33:43])
    IB write_data_pad_13 (.I(write_data[13]), .O(write_data_c_13));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(50[33:43])
    IB write_data_pad_12 (.I(write_data[12]), .O(write_data_c_12));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(50[33:43])
    IB write_data_pad_11 (.I(write_data[11]), .O(write_data_c_11));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(50[33:43])
    IB write_data_pad_10 (.I(write_data[10]), .O(write_data_c_10));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(50[33:43])
    IB write_data_pad_9 (.I(write_data[9]), .O(write_data_c_9));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(50[33:43])
    IB write_data_pad_8 (.I(write_data[8]), .O(write_data_c_8));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(50[33:43])
    IB write_data_pad_7 (.I(write_data[7]), .O(write_data_c_7));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(50[33:43])
    IB write_data_pad_6 (.I(write_data[6]), .O(write_data_c_6));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(50[33:43])
    IB write_data_pad_5 (.I(write_data[5]), .O(write_data_c_5));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(50[33:43])
    IB write_data_pad_4 (.I(write_data[4]), .O(write_data_c_4));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(50[33:43])
    IB write_data_pad_3 (.I(write_data[3]), .O(write_data_c_3));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(50[33:43])
    IB write_data_pad_2 (.I(write_data[2]), .O(write_data_c_2));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(50[33:43])
    IB write_data_pad_1 (.I(write_data[1]), .O(write_data_c_1));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(50[33:43])
    IB write_data_pad_0 (.I(write_data[0]), .O(write_data_c_0));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(50[33:43])
    FD1S3AX result_reg_i28 (.D(core_result[28]), .CK(clk_c), .Q(result_reg[28]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i28.GSR = "ENABLED";
    FD1S3AX result_reg_i29 (.D(core_result[29]), .CK(clk_c), .Q(result_reg[29]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i29.GSR = "ENABLED";
    FD1S3AX result_reg_i30 (.D(core_result[30]), .CK(clk_c), .Q(result_reg[30]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i30.GSR = "ENABLED";
    FD1S3AX result_reg_i31 (.D(core_result[31]), .CK(clk_c), .Q(result_reg[31]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i31.GSR = "ENABLED";
    FD1S3AX result_reg_i32 (.D(core_result[32]), .CK(clk_c), .Q(result_reg[32]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i32.GSR = "ENABLED";
    FD1S3AX result_reg_i33 (.D(core_result[33]), .CK(clk_c), .Q(result_reg[33]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i33.GSR = "ENABLED";
    FD1S3AX result_reg_i34 (.D(core_result[34]), .CK(clk_c), .Q(result_reg[34]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i34.GSR = "ENABLED";
    FD1S3AX result_reg_i35 (.D(core_result[35]), .CK(clk_c), .Q(result_reg[35]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i35.GSR = "ENABLED";
    FD1S3AX result_reg_i36 (.D(core_result[36]), .CK(clk_c), .Q(result_reg[36]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i36.GSR = "ENABLED";
    FD1S3AX result_reg_i37 (.D(core_result[37]), .CK(clk_c), .Q(result_reg[37]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i37.GSR = "ENABLED";
    FD1S3AX result_reg_i38 (.D(core_result[38]), .CK(clk_c), .Q(result_reg[38]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i38.GSR = "ENABLED";
    FD1S3AX result_reg_i39 (.D(core_result[39]), .CK(clk_c), .Q(result_reg[39]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i39.GSR = "ENABLED";
    FD1S3AX result_reg_i40 (.D(core_result[40]), .CK(clk_c), .Q(result_reg[40]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i40.GSR = "ENABLED";
    FD1S3AX result_reg_i41 (.D(core_result[41]), .CK(clk_c), .Q(result_reg[41]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i41.GSR = "ENABLED";
    FD1S3AX result_reg_i42 (.D(core_result[42]), .CK(clk_c), .Q(result_reg[42]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i42.GSR = "ENABLED";
    FD1S3AX result_reg_i43 (.D(core_result[43]), .CK(clk_c), .Q(result_reg[43]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i43.GSR = "ENABLED";
    FD1S3AX result_reg_i44 (.D(core_result[44]), .CK(clk_c), .Q(result_reg[44]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i44.GSR = "ENABLED";
    FD1S3AX result_reg_i45 (.D(core_result[45]), .CK(clk_c), .Q(result_reg[45]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i45.GSR = "ENABLED";
    FD1S3AX result_reg_i46 (.D(core_result[46]), .CK(clk_c), .Q(result_reg[46]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i46.GSR = "ENABLED";
    FD1S3AX result_reg_i47 (.D(core_result[47]), .CK(clk_c), .Q(result_reg[47]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i47.GSR = "ENABLED";
    FD1S3AX result_reg_i48 (.D(core_result[48]), .CK(clk_c), .Q(result_reg[48]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i48.GSR = "ENABLED";
    FD1S3AX result_reg_i49 (.D(core_result[49]), .CK(clk_c), .Q(result_reg[49]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i49.GSR = "ENABLED";
    FD1S3AX result_reg_i50 (.D(core_result[50]), .CK(clk_c), .Q(result_reg[50]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i50.GSR = "ENABLED";
    FD1S3AX result_reg_i51 (.D(core_result[51]), .CK(clk_c), .Q(result_reg[51]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i51.GSR = "ENABLED";
    FD1S3AX result_reg_i52 (.D(core_result[52]), .CK(clk_c), .Q(result_reg[52]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i52.GSR = "ENABLED";
    FD1S3AX result_reg_i53 (.D(core_result[53]), .CK(clk_c), .Q(result_reg[53]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i53.GSR = "ENABLED";
    FD1S3AX result_reg_i54 (.D(core_result[54]), .CK(clk_c), .Q(result_reg[54]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i54.GSR = "ENABLED";
    FD1S3AX result_reg_i55 (.D(core_result[55]), .CK(clk_c), .Q(result_reg[55]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i55.GSR = "ENABLED";
    FD1S3AX result_reg_i56 (.D(core_result[56]), .CK(clk_c), .Q(result_reg[56]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i56.GSR = "ENABLED";
    FD1S3AX result_reg_i57 (.D(core_result[57]), .CK(clk_c), .Q(result_reg[57]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i57.GSR = "ENABLED";
    FD1S3AX result_reg_i58 (.D(core_result[58]), .CK(clk_c), .Q(result_reg[58]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i58.GSR = "ENABLED";
    FD1S3AX result_reg_i59 (.D(core_result[59]), .CK(clk_c), .Q(result_reg[59]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i59.GSR = "ENABLED";
    FD1S3AX result_reg_i60 (.D(core_result[60]), .CK(clk_c), .Q(result_reg[60]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i60.GSR = "ENABLED";
    FD1S3AX result_reg_i61 (.D(core_result[61]), .CK(clk_c), .Q(result_reg[61]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i61.GSR = "ENABLED";
    FD1S3AX result_reg_i62 (.D(core_result[62]), .CK(clk_c), .Q(result_reg[62]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i62.GSR = "ENABLED";
    FD1S3AX result_reg_i63 (.D(core_result[63]), .CK(clk_c), .Q(result_reg[63]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i63.GSR = "ENABLED";
    FD1S3AX result_reg_i64 (.D(core_result[64]), .CK(clk_c), .Q(result_reg[64]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i64.GSR = "ENABLED";
    FD1S3AX result_reg_i65 (.D(core_result[65]), .CK(clk_c), .Q(result_reg[65]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i65.GSR = "ENABLED";
    FD1S3AX result_reg_i66 (.D(core_result[66]), .CK(clk_c), .Q(result_reg[66]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i66.GSR = "ENABLED";
    FD1S3AX result_reg_i67 (.D(core_result[67]), .CK(clk_c), .Q(result_reg[67]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i67.GSR = "ENABLED";
    FD1S3AX result_reg_i68 (.D(core_result[68]), .CK(clk_c), .Q(result_reg[68]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i68.GSR = "ENABLED";
    FD1S3AX result_reg_i69 (.D(core_result[69]), .CK(clk_c), .Q(result_reg[69]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i69.GSR = "ENABLED";
    FD1S3AX result_reg_i70 (.D(core_result[70]), .CK(clk_c), .Q(result_reg[70]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i70.GSR = "ENABLED";
    FD1S3AX result_reg_i71 (.D(core_result[71]), .CK(clk_c), .Q(result_reg[71]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i71.GSR = "ENABLED";
    FD1S3AX result_reg_i72 (.D(core_result[72]), .CK(clk_c), .Q(result_reg[72]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i72.GSR = "ENABLED";
    FD1S3AX result_reg_i73 (.D(core_result[73]), .CK(clk_c), .Q(result_reg[73]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i73.GSR = "ENABLED";
    FD1S3AX result_reg_i74 (.D(core_result[74]), .CK(clk_c), .Q(result_reg[74]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i74.GSR = "ENABLED";
    FD1S3AX result_reg_i75 (.D(core_result[75]), .CK(clk_c), .Q(result_reg[75]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i75.GSR = "ENABLED";
    FD1S3AX result_reg_i76 (.D(core_result[76]), .CK(clk_c), .Q(result_reg[76]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i76.GSR = "ENABLED";
    FD1S3AX result_reg_i77 (.D(core_result[77]), .CK(clk_c), .Q(result_reg[77]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i77.GSR = "ENABLED";
    FD1S3AX result_reg_i78 (.D(core_result[78]), .CK(clk_c), .Q(result_reg[78]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i78.GSR = "ENABLED";
    FD1S3AX result_reg_i79 (.D(core_result[79]), .CK(clk_c), .Q(result_reg[79]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i79.GSR = "ENABLED";
    FD1S3AX result_reg_i80 (.D(core_result[80]), .CK(clk_c), .Q(result_reg[80]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i80.GSR = "ENABLED";
    FD1S3AX result_reg_i81 (.D(core_result[81]), .CK(clk_c), .Q(result_reg[81]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i81.GSR = "ENABLED";
    FD1S3AX result_reg_i82 (.D(core_result[82]), .CK(clk_c), .Q(result_reg[82]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i82.GSR = "ENABLED";
    FD1S3AX result_reg_i83 (.D(core_result[83]), .CK(clk_c), .Q(result_reg[83]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i83.GSR = "ENABLED";
    FD1S3AX result_reg_i84 (.D(core_result[84]), .CK(clk_c), .Q(result_reg[84]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i84.GSR = "ENABLED";
    FD1S3AX result_reg_i85 (.D(core_result[85]), .CK(clk_c), .Q(result_reg[85]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i85.GSR = "ENABLED";
    FD1S3AX result_reg_i86 (.D(core_result[86]), .CK(clk_c), .Q(result_reg[86]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i86.GSR = "ENABLED";
    FD1S3AX result_reg_i87 (.D(core_result[87]), .CK(clk_c), .Q(result_reg[87]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i87.GSR = "ENABLED";
    FD1S3AX result_reg_i88 (.D(core_result[88]), .CK(clk_c), .Q(result_reg[88]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i88.GSR = "ENABLED";
    FD1S3AX result_reg_i89 (.D(core_result[89]), .CK(clk_c), .Q(result_reg[89]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i89.GSR = "ENABLED";
    FD1S3AX result_reg_i90 (.D(core_result[90]), .CK(clk_c), .Q(result_reg[90]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i90.GSR = "ENABLED";
    FD1S3AX result_reg_i91 (.D(core_result[91]), .CK(clk_c), .Q(result_reg[91]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i91.GSR = "ENABLED";
    FD1S3AX result_reg_i92 (.D(core_result[92]), .CK(clk_c), .Q(result_reg[92]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i92.GSR = "ENABLED";
    FD1S3AX result_reg_i93 (.D(core_result[93]), .CK(clk_c), .Q(result_reg[93]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i93.GSR = "ENABLED";
    FD1S3AX result_reg_i94 (.D(core_result[94]), .CK(clk_c), .Q(result_reg[94]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i94.GSR = "ENABLED";
    FD1S3AX result_reg_i95 (.D(core_result[95]), .CK(clk_c), .Q(result_reg[95]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i95.GSR = "ENABLED";
    FD1S3AX result_reg_i96 (.D(core_result[96]), .CK(clk_c), .Q(result_reg[96]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i96.GSR = "ENABLED";
    FD1S3AX result_reg_i97 (.D(core_result[97]), .CK(clk_c), .Q(result_reg[97]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i97.GSR = "ENABLED";
    FD1S3AX result_reg_i98 (.D(core_result[98]), .CK(clk_c), .Q(result_reg[98]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i98.GSR = "ENABLED";
    FD1S3AX result_reg_i99 (.D(core_result[99]), .CK(clk_c), .Q(result_reg[99]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i99.GSR = "ENABLED";
    FD1S3AX result_reg_i100 (.D(core_result[100]), .CK(clk_c), .Q(result_reg[100]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i100.GSR = "ENABLED";
    FD1S3AX result_reg_i101 (.D(core_result[101]), .CK(clk_c), .Q(result_reg[101]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i101.GSR = "ENABLED";
    FD1S3AX result_reg_i102 (.D(core_result[102]), .CK(clk_c), .Q(result_reg[102]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i102.GSR = "ENABLED";
    FD1S3AX result_reg_i103 (.D(core_result[103]), .CK(clk_c), .Q(result_reg[103]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i103.GSR = "ENABLED";
    FD1S3AX result_reg_i104 (.D(core_result[104]), .CK(clk_c), .Q(result_reg[104]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i104.GSR = "ENABLED";
    FD1S3AX result_reg_i105 (.D(core_result[105]), .CK(clk_c), .Q(result_reg[105]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i105.GSR = "ENABLED";
    FD1S3AX result_reg_i106 (.D(core_result[106]), .CK(clk_c), .Q(result_reg[106]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i106.GSR = "ENABLED";
    FD1S3AX result_reg_i107 (.D(core_result[107]), .CK(clk_c), .Q(result_reg[107]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i107.GSR = "ENABLED";
    FD1S3AX result_reg_i108 (.D(core_result[108]), .CK(clk_c), .Q(result_reg[108]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i108.GSR = "ENABLED";
    FD1S3AX result_reg_i109 (.D(core_result[109]), .CK(clk_c), .Q(result_reg[109]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i109.GSR = "ENABLED";
    FD1S3AX result_reg_i110 (.D(core_result[110]), .CK(clk_c), .Q(result_reg[110]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i110.GSR = "ENABLED";
    FD1S3AX result_reg_i111 (.D(core_result[111]), .CK(clk_c), .Q(result_reg[111]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i111.GSR = "ENABLED";
    FD1S3AX result_reg_i112 (.D(core_result[112]), .CK(clk_c), .Q(result_reg[112]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i112.GSR = "ENABLED";
    FD1S3AX result_reg_i113 (.D(core_result[113]), .CK(clk_c), .Q(result_reg[113]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i113.GSR = "ENABLED";
    FD1S3AX result_reg_i114 (.D(core_result[114]), .CK(clk_c), .Q(result_reg[114]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i114.GSR = "ENABLED";
    FD1S3AX result_reg_i115 (.D(core_result[115]), .CK(clk_c), .Q(result_reg[115]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i115.GSR = "ENABLED";
    FD1S3AX result_reg_i116 (.D(core_result[116]), .CK(clk_c), .Q(result_reg[116]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i116.GSR = "ENABLED";
    FD1S3AX result_reg_i117 (.D(core_result[117]), .CK(clk_c), .Q(result_reg[117]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i117.GSR = "ENABLED";
    FD1S3AX result_reg_i118 (.D(core_result[118]), .CK(clk_c), .Q(result_reg[118]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i118.GSR = "ENABLED";
    FD1S3AX result_reg_i119 (.D(core_result[119]), .CK(clk_c), .Q(result_reg[119]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i119.GSR = "ENABLED";
    FD1S3AX result_reg_i120 (.D(core_result[120]), .CK(clk_c), .Q(result_reg[120]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i120.GSR = "ENABLED";
    FD1S3AX result_reg_i121 (.D(core_result[121]), .CK(clk_c), .Q(result_reg[121]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i121.GSR = "ENABLED";
    FD1S3AX result_reg_i122 (.D(core_result[122]), .CK(clk_c), .Q(result_reg[122]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i122.GSR = "ENABLED";
    FD1S3AX result_reg_i123 (.D(core_result[123]), .CK(clk_c), .Q(result_reg[123]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i123.GSR = "ENABLED";
    FD1S3AX result_reg_i124 (.D(core_result[124]), .CK(clk_c), .Q(result_reg[124]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i124.GSR = "ENABLED";
    FD1S3AX result_reg_i125 (.D(core_result[125]), .CK(clk_c), .Q(result_reg[125]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i125.GSR = "ENABLED";
    FD1S3AX result_reg_i126 (.D(core_result[126]), .CK(clk_c), .Q(result_reg[126]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i126.GSR = "ENABLED";
    FD1S3AX result_reg_i127 (.D(core_result[127]), .CK(clk_c), .Q(result_reg[127]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam result_reg_i127.GSR = "ENABLED";
    PFUMX i29050 (.BLUT(n34001), .ALUT(n34002), .C0(address_c_0), .Z(n34003));
    FD1P3AX key_reg_7___i2 (.D(write_data_c_1), .SP(clk_c_enable_163), .CK(clk_c), 
            .Q(\key_reg[7] [1]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i2.GSR = "ENABLED";
    FD1P3AX key_reg_7___i3 (.D(write_data_c_2), .SP(clk_c_enable_163), .CK(clk_c), 
            .Q(\key_reg[7] [2]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i3.GSR = "ENABLED";
    FD1P3AX key_reg_7___i4 (.D(write_data_c_3), .SP(clk_c_enable_163), .CK(clk_c), 
            .Q(\key_reg[7] [3]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i4.GSR = "ENABLED";
    FD1P3AX key_reg_7___i5 (.D(write_data_c_4), .SP(clk_c_enable_163), .CK(clk_c), 
            .Q(\key_reg[7] [4]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i5.GSR = "ENABLED";
    FD1P3AX key_reg_7___i6 (.D(write_data_c_5), .SP(clk_c_enable_163), .CK(clk_c), 
            .Q(\key_reg[7] [5]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i6.GSR = "ENABLED";
    FD1P3AX key_reg_7___i7 (.D(write_data_c_6), .SP(clk_c_enable_163), .CK(clk_c), 
            .Q(\key_reg[7] [6]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i7.GSR = "ENABLED";
    FD1P3AX key_reg_7___i8 (.D(write_data_c_7), .SP(clk_c_enable_163), .CK(clk_c), 
            .Q(\key_reg[7] [7]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i8.GSR = "ENABLED";
    FD1P3AX key_reg_7___i9 (.D(write_data_c_8), .SP(clk_c_enable_163), .CK(clk_c), 
            .Q(\key_reg[7] [8]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i9.GSR = "ENABLED";
    FD1P3AX key_reg_7___i10 (.D(write_data_c_9), .SP(clk_c_enable_163), 
            .CK(clk_c), .Q(\key_reg[7] [9]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i10.GSR = "ENABLED";
    FD1P3AX key_reg_7___i11 (.D(write_data_c_10), .SP(clk_c_enable_163), 
            .CK(clk_c), .Q(\key_reg[7] [10]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i11.GSR = "ENABLED";
    FD1P3AX key_reg_7___i12 (.D(write_data_c_11), .SP(clk_c_enable_163), 
            .CK(clk_c), .Q(\key_reg[7] [11]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i12.GSR = "ENABLED";
    FD1P3AX key_reg_7___i13 (.D(write_data_c_12), .SP(clk_c_enable_163), 
            .CK(clk_c), .Q(\key_reg[7] [12]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i13.GSR = "ENABLED";
    FD1P3AX key_reg_7___i14 (.D(write_data_c_13), .SP(clk_c_enable_163), 
            .CK(clk_c), .Q(\key_reg[7] [13]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i14.GSR = "ENABLED";
    FD1P3AX key_reg_7___i15 (.D(write_data_c_14), .SP(clk_c_enable_163), 
            .CK(clk_c), .Q(\key_reg[7] [14]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i15.GSR = "ENABLED";
    FD1P3AX key_reg_7___i16 (.D(write_data_c_15), .SP(clk_c_enable_163), 
            .CK(clk_c), .Q(\key_reg[7] [15]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i16.GSR = "ENABLED";
    FD1P3AX key_reg_7___i17 (.D(write_data_c_16), .SP(clk_c_enable_163), 
            .CK(clk_c), .Q(\key_reg[7] [16]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i17.GSR = "ENABLED";
    FD1P3AX key_reg_7___i18 (.D(write_data_c_17), .SP(clk_c_enable_163), 
            .CK(clk_c), .Q(\key_reg[7] [17]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i18.GSR = "ENABLED";
    FD1P3AX key_reg_7___i19 (.D(write_data_c_18), .SP(clk_c_enable_163), 
            .CK(clk_c), .Q(\key_reg[7] [18]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i19.GSR = "ENABLED";
    FD1P3AX key_reg_7___i20 (.D(write_data_c_19), .SP(clk_c_enable_163), 
            .CK(clk_c), .Q(\key_reg[7] [19]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i20.GSR = "ENABLED";
    FD1P3AX key_reg_7___i21 (.D(write_data_c_20), .SP(clk_c_enable_163), 
            .CK(clk_c), .Q(\key_reg[7] [20]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i21.GSR = "ENABLED";
    FD1P3AX key_reg_7___i22 (.D(write_data_c_21), .SP(clk_c_enable_163), 
            .CK(clk_c), .Q(\key_reg[7] [21]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i22.GSR = "ENABLED";
    FD1P3AX key_reg_7___i23 (.D(write_data_c_22), .SP(clk_c_enable_163), 
            .CK(clk_c), .Q(\key_reg[7] [22]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i23.GSR = "ENABLED";
    FD1P3AX key_reg_7___i24 (.D(write_data_c_23), .SP(clk_c_enable_163), 
            .CK(clk_c), .Q(\key_reg[7] [23]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i24.GSR = "ENABLED";
    FD1P3AX key_reg_7___i25 (.D(write_data_c_24), .SP(clk_c_enable_163), 
            .CK(clk_c), .Q(\key_reg[7] [24]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i25.GSR = "ENABLED";
    FD1P3AX key_reg_7___i26 (.D(write_data_c_25), .SP(clk_c_enable_163), 
            .CK(clk_c), .Q(\key_reg[7] [25]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i26.GSR = "ENABLED";
    FD1P3AX key_reg_7___i27 (.D(write_data_c_26), .SP(clk_c_enable_163), 
            .CK(clk_c), .Q(\key_reg[7] [26]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i27.GSR = "ENABLED";
    FD1P3AX key_reg_7___i28 (.D(write_data_c_27), .SP(clk_c_enable_163), 
            .CK(clk_c), .Q(\key_reg[7] [27]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i28.GSR = "ENABLED";
    FD1P3AX key_reg_7___i29 (.D(write_data_c_28), .SP(clk_c_enable_163), 
            .CK(clk_c), .Q(\key_reg[7] [28]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i29.GSR = "ENABLED";
    FD1P3AX key_reg_7___i30 (.D(write_data_c_29), .SP(clk_c_enable_163), 
            .CK(clk_c), .Q(\key_reg[7] [29]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i30.GSR = "ENABLED";
    FD1P3AX key_reg_7___i31 (.D(write_data_c_30), .SP(clk_c_enable_163), 
            .CK(clk_c), .Q(\key_reg[7] [30]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i31.GSR = "ENABLED";
    FD1P3AX key_reg_7___i32 (.D(write_data_c_31), .SP(clk_c_enable_163), 
            .CK(clk_c), .Q(\key_reg[7] [31]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i32.GSR = "ENABLED";
    FD1P3AX key_reg_7___i33 (.D(write_data_c_0), .SP(clk_c_enable_195), 
            .CK(clk_c), .Q(\key_reg[6] [0]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i33.GSR = "ENABLED";
    FD1P3AX key_reg_7___i34 (.D(write_data_c_1), .SP(clk_c_enable_195), 
            .CK(clk_c), .Q(\key_reg[6] [1]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i34.GSR = "ENABLED";
    FD1P3AX key_reg_7___i35 (.D(write_data_c_2), .SP(clk_c_enable_195), 
            .CK(clk_c), .Q(\key_reg[6] [2]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i35.GSR = "ENABLED";
    FD1P3AX key_reg_7___i36 (.D(write_data_c_3), .SP(clk_c_enable_195), 
            .CK(clk_c), .Q(\key_reg[6] [3]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i36.GSR = "ENABLED";
    FD1P3AX key_reg_7___i37 (.D(write_data_c_4), .SP(clk_c_enable_195), 
            .CK(clk_c), .Q(\key_reg[6] [4]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i37.GSR = "ENABLED";
    FD1P3AX key_reg_7___i38 (.D(write_data_c_5), .SP(clk_c_enable_195), 
            .CK(clk_c), .Q(\key_reg[6] [5]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i38.GSR = "ENABLED";
    FD1P3AX key_reg_7___i39 (.D(write_data_c_6), .SP(clk_c_enable_195), 
            .CK(clk_c), .Q(\key_reg[6] [6]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i39.GSR = "ENABLED";
    FD1P3AX key_reg_7___i40 (.D(write_data_c_7), .SP(clk_c_enable_195), 
            .CK(clk_c), .Q(\key_reg[6] [7]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i40.GSR = "ENABLED";
    FD1P3AX key_reg_7___i41 (.D(write_data_c_8), .SP(clk_c_enable_195), 
            .CK(clk_c), .Q(\key_reg[6] [8]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i41.GSR = "ENABLED";
    FD1P3AX key_reg_7___i42 (.D(write_data_c_9), .SP(clk_c_enable_195), 
            .CK(clk_c), .Q(\key_reg[6] [9]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i42.GSR = "ENABLED";
    FD1P3AX key_reg_7___i43 (.D(write_data_c_10), .SP(clk_c_enable_195), 
            .CK(clk_c), .Q(\key_reg[6] [10]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i43.GSR = "ENABLED";
    FD1P3AX key_reg_7___i44 (.D(write_data_c_11), .SP(clk_c_enable_195), 
            .CK(clk_c), .Q(\key_reg[6] [11]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i44.GSR = "ENABLED";
    FD1P3AX key_reg_7___i45 (.D(write_data_c_12), .SP(clk_c_enable_195), 
            .CK(clk_c), .Q(\key_reg[6] [12]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i45.GSR = "ENABLED";
    FD1P3AX key_reg_7___i46 (.D(write_data_c_13), .SP(clk_c_enable_195), 
            .CK(clk_c), .Q(\key_reg[6] [13]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i46.GSR = "ENABLED";
    FD1P3AX key_reg_7___i47 (.D(write_data_c_14), .SP(clk_c_enable_195), 
            .CK(clk_c), .Q(\key_reg[6] [14]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i47.GSR = "ENABLED";
    FD1P3AX key_reg_7___i48 (.D(write_data_c_15), .SP(clk_c_enable_195), 
            .CK(clk_c), .Q(\key_reg[6] [15]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i48.GSR = "ENABLED";
    FD1P3AX key_reg_7___i49 (.D(write_data_c_16), .SP(clk_c_enable_195), 
            .CK(clk_c), .Q(\key_reg[6] [16]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i49.GSR = "ENABLED";
    FD1P3AX key_reg_7___i50 (.D(write_data_c_17), .SP(clk_c_enable_195), 
            .CK(clk_c), .Q(\key_reg[6] [17]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i50.GSR = "ENABLED";
    FD1P3AX key_reg_7___i51 (.D(write_data_c_18), .SP(clk_c_enable_195), 
            .CK(clk_c), .Q(\key_reg[6] [18]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i51.GSR = "ENABLED";
    FD1P3AX key_reg_7___i52 (.D(write_data_c_19), .SP(clk_c_enable_195), 
            .CK(clk_c), .Q(\key_reg[6] [19]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i52.GSR = "ENABLED";
    FD1P3AX key_reg_7___i53 (.D(write_data_c_20), .SP(clk_c_enable_195), 
            .CK(clk_c), .Q(\key_reg[6] [20]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i53.GSR = "ENABLED";
    FD1P3AX key_reg_7___i54 (.D(write_data_c_21), .SP(clk_c_enable_195), 
            .CK(clk_c), .Q(\key_reg[6] [21]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i54.GSR = "ENABLED";
    FD1P3AX key_reg_7___i55 (.D(write_data_c_22), .SP(clk_c_enable_195), 
            .CK(clk_c), .Q(\key_reg[6] [22]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i55.GSR = "ENABLED";
    FD1P3AX key_reg_7___i56 (.D(write_data_c_23), .SP(clk_c_enable_195), 
            .CK(clk_c), .Q(\key_reg[6] [23]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i56.GSR = "ENABLED";
    FD1P3AX key_reg_7___i57 (.D(write_data_c_24), .SP(clk_c_enable_195), 
            .CK(clk_c), .Q(\key_reg[6] [24]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i57.GSR = "ENABLED";
    FD1P3AX key_reg_7___i58 (.D(write_data_c_25), .SP(clk_c_enable_195), 
            .CK(clk_c), .Q(\key_reg[6] [25]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i58.GSR = "ENABLED";
    FD1P3AX key_reg_7___i59 (.D(write_data_c_26), .SP(clk_c_enable_195), 
            .CK(clk_c), .Q(\key_reg[6] [26]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i59.GSR = "ENABLED";
    FD1P3AX key_reg_7___i60 (.D(write_data_c_27), .SP(clk_c_enable_195), 
            .CK(clk_c), .Q(\key_reg[6] [27]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i60.GSR = "ENABLED";
    FD1P3AX key_reg_7___i61 (.D(write_data_c_28), .SP(clk_c_enable_195), 
            .CK(clk_c), .Q(\key_reg[6] [28]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i61.GSR = "ENABLED";
    FD1P3AX key_reg_7___i62 (.D(write_data_c_29), .SP(clk_c_enable_195), 
            .CK(clk_c), .Q(\key_reg[6] [29]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i62.GSR = "ENABLED";
    FD1P3AX key_reg_7___i63 (.D(write_data_c_30), .SP(clk_c_enable_195), 
            .CK(clk_c), .Q(\key_reg[6] [30]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i63.GSR = "ENABLED";
    FD1P3AX key_reg_7___i64 (.D(write_data_c_31), .SP(clk_c_enable_195), 
            .CK(clk_c), .Q(\key_reg[6] [31]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i64.GSR = "ENABLED";
    FD1P3AX key_reg_7___i65 (.D(write_data_c_0), .SP(clk_c_enable_227), 
            .CK(clk_c), .Q(\key_reg[5] [0]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i65.GSR = "ENABLED";
    FD1P3AX key_reg_7___i66 (.D(write_data_c_1), .SP(clk_c_enable_227), 
            .CK(clk_c), .Q(\key_reg[5] [1]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i66.GSR = "ENABLED";
    FD1P3AX key_reg_7___i67 (.D(write_data_c_2), .SP(clk_c_enable_227), 
            .CK(clk_c), .Q(\key_reg[5] [2]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i67.GSR = "ENABLED";
    FD1P3AX key_reg_7___i68 (.D(write_data_c_3), .SP(clk_c_enable_227), 
            .CK(clk_c), .Q(\key_reg[5] [3]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i68.GSR = "ENABLED";
    FD1P3AX key_reg_7___i69 (.D(write_data_c_4), .SP(clk_c_enable_227), 
            .CK(clk_c), .Q(\key_reg[5] [4]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i69.GSR = "ENABLED";
    FD1P3AX key_reg_7___i70 (.D(write_data_c_5), .SP(clk_c_enable_227), 
            .CK(clk_c), .Q(\key_reg[5] [5]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i70.GSR = "ENABLED";
    FD1P3AX key_reg_7___i71 (.D(write_data_c_6), .SP(clk_c_enable_227), 
            .CK(clk_c), .Q(\key_reg[5] [6]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i71.GSR = "ENABLED";
    FD1P3AX key_reg_7___i72 (.D(write_data_c_7), .SP(clk_c_enable_227), 
            .CK(clk_c), .Q(\key_reg[5] [7]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i72.GSR = "ENABLED";
    FD1P3AX key_reg_7___i73 (.D(write_data_c_8), .SP(clk_c_enable_227), 
            .CK(clk_c), .Q(\key_reg[5] [8]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i73.GSR = "ENABLED";
    FD1P3AX key_reg_7___i74 (.D(write_data_c_9), .SP(clk_c_enable_227), 
            .CK(clk_c), .Q(\key_reg[5] [9]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i74.GSR = "ENABLED";
    FD1P3AX key_reg_7___i75 (.D(write_data_c_10), .SP(clk_c_enable_227), 
            .CK(clk_c), .Q(\key_reg[5] [10]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i75.GSR = "ENABLED";
    FD1P3AX key_reg_7___i76 (.D(write_data_c_11), .SP(clk_c_enable_227), 
            .CK(clk_c), .Q(\key_reg[5] [11]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i76.GSR = "ENABLED";
    FD1P3AX key_reg_7___i77 (.D(write_data_c_12), .SP(clk_c_enable_227), 
            .CK(clk_c), .Q(\key_reg[5] [12]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i77.GSR = "ENABLED";
    FD1P3AX key_reg_7___i78 (.D(write_data_c_13), .SP(clk_c_enable_227), 
            .CK(clk_c), .Q(\key_reg[5] [13]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i78.GSR = "ENABLED";
    FD1P3AX key_reg_7___i79 (.D(write_data_c_14), .SP(clk_c_enable_227), 
            .CK(clk_c), .Q(\key_reg[5] [14]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i79.GSR = "ENABLED";
    FD1P3AX key_reg_7___i80 (.D(write_data_c_15), .SP(clk_c_enable_227), 
            .CK(clk_c), .Q(\key_reg[5] [15]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i80.GSR = "ENABLED";
    FD1P3AX key_reg_7___i81 (.D(write_data_c_16), .SP(clk_c_enable_227), 
            .CK(clk_c), .Q(\key_reg[5] [16]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i81.GSR = "ENABLED";
    FD1P3AX key_reg_7___i82 (.D(write_data_c_17), .SP(clk_c_enable_227), 
            .CK(clk_c), .Q(\key_reg[5] [17]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i82.GSR = "ENABLED";
    FD1P3AX key_reg_7___i83 (.D(write_data_c_18), .SP(clk_c_enable_227), 
            .CK(clk_c), .Q(\key_reg[5] [18]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i83.GSR = "ENABLED";
    FD1P3AX key_reg_7___i84 (.D(write_data_c_19), .SP(clk_c_enable_227), 
            .CK(clk_c), .Q(\key_reg[5] [19]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i84.GSR = "ENABLED";
    FD1P3AX key_reg_7___i85 (.D(write_data_c_20), .SP(clk_c_enable_227), 
            .CK(clk_c), .Q(\key_reg[5] [20]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i85.GSR = "ENABLED";
    FD1P3AX key_reg_7___i86 (.D(write_data_c_21), .SP(clk_c_enable_227), 
            .CK(clk_c), .Q(\key_reg[5] [21]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i86.GSR = "ENABLED";
    FD1P3AX key_reg_7___i87 (.D(write_data_c_22), .SP(clk_c_enable_227), 
            .CK(clk_c), .Q(\key_reg[5] [22]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i87.GSR = "ENABLED";
    FD1P3AX key_reg_7___i88 (.D(write_data_c_23), .SP(clk_c_enable_227), 
            .CK(clk_c), .Q(\key_reg[5] [23]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i88.GSR = "ENABLED";
    FD1P3AX key_reg_7___i89 (.D(write_data_c_24), .SP(clk_c_enable_227), 
            .CK(clk_c), .Q(\key_reg[5] [24]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i89.GSR = "ENABLED";
    FD1P3AX key_reg_7___i90 (.D(write_data_c_25), .SP(clk_c_enable_227), 
            .CK(clk_c), .Q(\key_reg[5] [25]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i90.GSR = "ENABLED";
    FD1P3AX key_reg_7___i91 (.D(write_data_c_26), .SP(clk_c_enable_227), 
            .CK(clk_c), .Q(\key_reg[5] [26]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i91.GSR = "ENABLED";
    FD1P3AX key_reg_7___i92 (.D(write_data_c_27), .SP(clk_c_enable_227), 
            .CK(clk_c), .Q(\key_reg[5] [27]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i92.GSR = "ENABLED";
    FD1P3AX key_reg_7___i93 (.D(write_data_c_28), .SP(clk_c_enable_227), 
            .CK(clk_c), .Q(\key_reg[5] [28]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i93.GSR = "ENABLED";
    FD1P3AX key_reg_7___i94 (.D(write_data_c_29), .SP(clk_c_enable_227), 
            .CK(clk_c), .Q(\key_reg[5] [29]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i94.GSR = "ENABLED";
    FD1P3AX key_reg_7___i95 (.D(write_data_c_30), .SP(clk_c_enable_227), 
            .CK(clk_c), .Q(\key_reg[5] [30]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i95.GSR = "ENABLED";
    FD1P3AX key_reg_7___i96 (.D(write_data_c_31), .SP(clk_c_enable_227), 
            .CK(clk_c), .Q(\key_reg[5] [31]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i96.GSR = "ENABLED";
    FD1P3AX key_reg_7___i97 (.D(write_data_c_0), .SP(clk_c_enable_259), 
            .CK(clk_c), .Q(\key_reg[4] [0]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i97.GSR = "ENABLED";
    FD1P3AX key_reg_7___i98 (.D(write_data_c_1), .SP(clk_c_enable_259), 
            .CK(clk_c), .Q(\key_reg[4] [1]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i98.GSR = "ENABLED";
    FD1P3AX key_reg_7___i99 (.D(write_data_c_2), .SP(clk_c_enable_259), 
            .CK(clk_c), .Q(\key_reg[4] [2]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i99.GSR = "ENABLED";
    FD1P3AX key_reg_7___i100 (.D(write_data_c_3), .SP(clk_c_enable_259), 
            .CK(clk_c), .Q(\key_reg[4] [3]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i100.GSR = "ENABLED";
    FD1P3AX key_reg_7___i101 (.D(write_data_c_4), .SP(clk_c_enable_259), 
            .CK(clk_c), .Q(\key_reg[4] [4]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i101.GSR = "ENABLED";
    FD1P3AX key_reg_7___i102 (.D(write_data_c_5), .SP(clk_c_enable_259), 
            .CK(clk_c), .Q(\key_reg[4] [5]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i102.GSR = "ENABLED";
    FD1P3AX key_reg_7___i103 (.D(write_data_c_6), .SP(clk_c_enable_259), 
            .CK(clk_c), .Q(\key_reg[4] [6]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i103.GSR = "ENABLED";
    FD1P3AX key_reg_7___i104 (.D(write_data_c_7), .SP(clk_c_enable_259), 
            .CK(clk_c), .Q(\key_reg[4] [7]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i104.GSR = "ENABLED";
    FD1P3AX key_reg_7___i105 (.D(write_data_c_8), .SP(clk_c_enable_259), 
            .CK(clk_c), .Q(\key_reg[4] [8]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i105.GSR = "ENABLED";
    FD1P3AX key_reg_7___i106 (.D(write_data_c_9), .SP(clk_c_enable_259), 
            .CK(clk_c), .Q(\key_reg[4] [9]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i106.GSR = "ENABLED";
    FD1P3AX key_reg_7___i107 (.D(write_data_c_10), .SP(clk_c_enable_259), 
            .CK(clk_c), .Q(\key_reg[4] [10]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i107.GSR = "ENABLED";
    FD1P3AX key_reg_7___i108 (.D(write_data_c_11), .SP(clk_c_enable_259), 
            .CK(clk_c), .Q(\key_reg[4] [11]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i108.GSR = "ENABLED";
    FD1P3AX key_reg_7___i109 (.D(write_data_c_12), .SP(clk_c_enable_259), 
            .CK(clk_c), .Q(\key_reg[4] [12]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i109.GSR = "ENABLED";
    FD1P3AX key_reg_7___i110 (.D(write_data_c_13), .SP(clk_c_enable_259), 
            .CK(clk_c), .Q(\key_reg[4] [13]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i110.GSR = "ENABLED";
    FD1P3AX key_reg_7___i111 (.D(write_data_c_14), .SP(clk_c_enable_259), 
            .CK(clk_c), .Q(\key_reg[4] [14]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i111.GSR = "ENABLED";
    FD1P3AX key_reg_7___i112 (.D(write_data_c_15), .SP(clk_c_enable_259), 
            .CK(clk_c), .Q(\key_reg[4] [15]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i112.GSR = "ENABLED";
    FD1P3AX key_reg_7___i113 (.D(write_data_c_16), .SP(clk_c_enable_259), 
            .CK(clk_c), .Q(\key_reg[4] [16]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i113.GSR = "ENABLED";
    FD1P3AX key_reg_7___i114 (.D(write_data_c_17), .SP(clk_c_enable_259), 
            .CK(clk_c), .Q(\key_reg[4] [17]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i114.GSR = "ENABLED";
    FD1P3AX key_reg_7___i115 (.D(write_data_c_18), .SP(clk_c_enable_259), 
            .CK(clk_c), .Q(\key_reg[4] [18]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i115.GSR = "ENABLED";
    FD1P3AX key_reg_7___i116 (.D(write_data_c_19), .SP(clk_c_enable_259), 
            .CK(clk_c), .Q(\key_reg[4] [19]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i116.GSR = "ENABLED";
    FD1P3AX key_reg_7___i117 (.D(write_data_c_20), .SP(clk_c_enable_259), 
            .CK(clk_c), .Q(\key_reg[4] [20]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i117.GSR = "ENABLED";
    FD1P3AX key_reg_7___i118 (.D(write_data_c_21), .SP(clk_c_enable_259), 
            .CK(clk_c), .Q(\key_reg[4] [21]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i118.GSR = "ENABLED";
    FD1P3AX key_reg_7___i119 (.D(write_data_c_22), .SP(clk_c_enable_259), 
            .CK(clk_c), .Q(\key_reg[4] [22]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i119.GSR = "ENABLED";
    FD1P3AX key_reg_7___i120 (.D(write_data_c_23), .SP(clk_c_enable_259), 
            .CK(clk_c), .Q(\key_reg[4] [23]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i120.GSR = "ENABLED";
    FD1P3AX key_reg_7___i121 (.D(write_data_c_24), .SP(clk_c_enable_259), 
            .CK(clk_c), .Q(\key_reg[4] [24]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i121.GSR = "ENABLED";
    FD1P3AX key_reg_7___i122 (.D(write_data_c_25), .SP(clk_c_enable_259), 
            .CK(clk_c), .Q(\key_reg[4] [25]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i122.GSR = "ENABLED";
    FD1P3AX key_reg_7___i123 (.D(write_data_c_26), .SP(clk_c_enable_259), 
            .CK(clk_c), .Q(\key_reg[4] [26]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i123.GSR = "ENABLED";
    FD1P3AX key_reg_7___i124 (.D(write_data_c_27), .SP(clk_c_enable_259), 
            .CK(clk_c), .Q(\key_reg[4] [27]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i124.GSR = "ENABLED";
    FD1P3AX key_reg_7___i125 (.D(write_data_c_28), .SP(clk_c_enable_259), 
            .CK(clk_c), .Q(\key_reg[4] [28]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i125.GSR = "ENABLED";
    FD1P3AX key_reg_7___i126 (.D(write_data_c_29), .SP(clk_c_enable_259), 
            .CK(clk_c), .Q(\key_reg[4] [29]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i126.GSR = "ENABLED";
    FD1P3AX key_reg_7___i127 (.D(write_data_c_30), .SP(clk_c_enable_259), 
            .CK(clk_c), .Q(\key_reg[4] [30]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i127.GSR = "ENABLED";
    FD1P3AX key_reg_7___i128 (.D(write_data_c_31), .SP(clk_c_enable_259), 
            .CK(clk_c), .Q(\key_reg[4] [31]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i128.GSR = "ENABLED";
    FD1P3AX key_reg_7___i129 (.D(write_data_c_0), .SP(clk_c_enable_291), 
            .CK(clk_c), .Q(\key_reg[3] [0]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i129.GSR = "ENABLED";
    FD1P3AX key_reg_7___i130 (.D(write_data_c_1), .SP(clk_c_enable_291), 
            .CK(clk_c), .Q(\key_reg[3] [1]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i130.GSR = "ENABLED";
    FD1P3AX key_reg_7___i131 (.D(write_data_c_2), .SP(clk_c_enable_291), 
            .CK(clk_c), .Q(\key_reg[3] [2]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i131.GSR = "ENABLED";
    FD1P3AX key_reg_7___i132 (.D(write_data_c_3), .SP(clk_c_enable_291), 
            .CK(clk_c), .Q(\key_reg[3] [3]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i132.GSR = "ENABLED";
    FD1P3AX key_reg_7___i133 (.D(write_data_c_4), .SP(clk_c_enable_291), 
            .CK(clk_c), .Q(\key_reg[3] [4]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i133.GSR = "ENABLED";
    FD1P3AX key_reg_7___i134 (.D(write_data_c_5), .SP(clk_c_enable_291), 
            .CK(clk_c), .Q(\key_reg[3] [5]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i134.GSR = "ENABLED";
    FD1P3AX key_reg_7___i135 (.D(write_data_c_6), .SP(clk_c_enable_291), 
            .CK(clk_c), .Q(\key_reg[3] [6]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i135.GSR = "ENABLED";
    FD1P3AX key_reg_7___i136 (.D(write_data_c_7), .SP(clk_c_enable_291), 
            .CK(clk_c), .Q(\key_reg[3] [7]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i136.GSR = "ENABLED";
    FD1P3AX key_reg_7___i137 (.D(write_data_c_8), .SP(clk_c_enable_291), 
            .CK(clk_c), .Q(\key_reg[3] [8]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i137.GSR = "ENABLED";
    FD1P3AX key_reg_7___i138 (.D(write_data_c_9), .SP(clk_c_enable_291), 
            .CK(clk_c), .Q(\key_reg[3] [9]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i138.GSR = "ENABLED";
    FD1P3AX key_reg_7___i139 (.D(write_data_c_10), .SP(clk_c_enable_291), 
            .CK(clk_c), .Q(\key_reg[3] [10]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i139.GSR = "ENABLED";
    FD1P3AX key_reg_7___i140 (.D(write_data_c_11), .SP(clk_c_enable_291), 
            .CK(clk_c), .Q(\key_reg[3] [11]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i140.GSR = "ENABLED";
    FD1P3AX key_reg_7___i141 (.D(write_data_c_12), .SP(clk_c_enable_291), 
            .CK(clk_c), .Q(\key_reg[3] [12]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i141.GSR = "ENABLED";
    FD1P3AX key_reg_7___i142 (.D(write_data_c_13), .SP(clk_c_enable_291), 
            .CK(clk_c), .Q(\key_reg[3] [13]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i142.GSR = "ENABLED";
    FD1P3AX key_reg_7___i143 (.D(write_data_c_14), .SP(clk_c_enable_291), 
            .CK(clk_c), .Q(\key_reg[3] [14]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i143.GSR = "ENABLED";
    FD1P3AX key_reg_7___i144 (.D(write_data_c_15), .SP(clk_c_enable_291), 
            .CK(clk_c), .Q(\key_reg[3] [15]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i144.GSR = "ENABLED";
    FD1P3AX key_reg_7___i145 (.D(write_data_c_16), .SP(clk_c_enable_291), 
            .CK(clk_c), .Q(\key_reg[3] [16]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i145.GSR = "ENABLED";
    FD1P3AX key_reg_7___i146 (.D(write_data_c_17), .SP(clk_c_enable_291), 
            .CK(clk_c), .Q(\key_reg[3] [17]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i146.GSR = "ENABLED";
    FD1P3AX key_reg_7___i147 (.D(write_data_c_18), .SP(clk_c_enable_291), 
            .CK(clk_c), .Q(\key_reg[3] [18]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i147.GSR = "ENABLED";
    FD1P3AX key_reg_7___i148 (.D(write_data_c_19), .SP(clk_c_enable_291), 
            .CK(clk_c), .Q(\key_reg[3] [19]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i148.GSR = "ENABLED";
    FD1P3AX key_reg_7___i149 (.D(write_data_c_20), .SP(clk_c_enable_291), 
            .CK(clk_c), .Q(\key_reg[3] [20]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i149.GSR = "ENABLED";
    FD1P3AX key_reg_7___i150 (.D(write_data_c_21), .SP(clk_c_enable_291), 
            .CK(clk_c), .Q(\key_reg[3] [21]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i150.GSR = "ENABLED";
    FD1P3AX key_reg_7___i151 (.D(write_data_c_22), .SP(clk_c_enable_291), 
            .CK(clk_c), .Q(\key_reg[3] [22]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i151.GSR = "ENABLED";
    FD1P3AX key_reg_7___i152 (.D(write_data_c_23), .SP(clk_c_enable_291), 
            .CK(clk_c), .Q(\key_reg[3] [23]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i152.GSR = "ENABLED";
    FD1P3AX key_reg_7___i153 (.D(write_data_c_24), .SP(clk_c_enable_291), 
            .CK(clk_c), .Q(\key_reg[3] [24]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i153.GSR = "ENABLED";
    FD1P3AX key_reg_7___i154 (.D(write_data_c_25), .SP(clk_c_enable_291), 
            .CK(clk_c), .Q(\key_reg[3] [25]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i154.GSR = "ENABLED";
    FD1P3AX key_reg_7___i155 (.D(write_data_c_26), .SP(clk_c_enable_291), 
            .CK(clk_c), .Q(\key_reg[3] [26]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i155.GSR = "ENABLED";
    FD1P3AX key_reg_7___i156 (.D(write_data_c_27), .SP(clk_c_enable_291), 
            .CK(clk_c), .Q(\key_reg[3] [27]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i156.GSR = "ENABLED";
    FD1P3AX key_reg_7___i157 (.D(write_data_c_28), .SP(clk_c_enable_291), 
            .CK(clk_c), .Q(\key_reg[3] [28]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i157.GSR = "ENABLED";
    FD1P3AX key_reg_7___i158 (.D(write_data_c_29), .SP(clk_c_enable_291), 
            .CK(clk_c), .Q(\key_reg[3] [29]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i158.GSR = "ENABLED";
    FD1P3AX key_reg_7___i159 (.D(write_data_c_30), .SP(clk_c_enable_291), 
            .CK(clk_c), .Q(\key_reg[3] [30]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i159.GSR = "ENABLED";
    FD1P3AX key_reg_7___i160 (.D(write_data_c_31), .SP(clk_c_enable_291), 
            .CK(clk_c), .Q(\key_reg[3] [31]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i160.GSR = "ENABLED";
    FD1P3AX key_reg_7___i161 (.D(write_data_c_0), .SP(clk_c_enable_323), 
            .CK(clk_c), .Q(\key_reg[2] [0]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i161.GSR = "ENABLED";
    FD1P3AX key_reg_7___i162 (.D(write_data_c_1), .SP(clk_c_enable_323), 
            .CK(clk_c), .Q(\key_reg[2] [1]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i162.GSR = "ENABLED";
    FD1P3AX key_reg_7___i163 (.D(write_data_c_2), .SP(clk_c_enable_323), 
            .CK(clk_c), .Q(\key_reg[2] [2]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i163.GSR = "ENABLED";
    FD1P3AX key_reg_7___i164 (.D(write_data_c_3), .SP(clk_c_enable_323), 
            .CK(clk_c), .Q(\key_reg[2] [3]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i164.GSR = "ENABLED";
    FD1P3AX key_reg_7___i165 (.D(write_data_c_4), .SP(clk_c_enable_323), 
            .CK(clk_c), .Q(\key_reg[2] [4]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i165.GSR = "ENABLED";
    FD1P3AX key_reg_7___i166 (.D(write_data_c_5), .SP(clk_c_enable_323), 
            .CK(clk_c), .Q(\key_reg[2] [5]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i166.GSR = "ENABLED";
    FD1P3AX key_reg_7___i167 (.D(write_data_c_6), .SP(clk_c_enable_323), 
            .CK(clk_c), .Q(\key_reg[2] [6]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i167.GSR = "ENABLED";
    FD1P3AX key_reg_7___i168 (.D(write_data_c_7), .SP(clk_c_enable_323), 
            .CK(clk_c), .Q(\key_reg[2] [7]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i168.GSR = "ENABLED";
    FD1P3AX key_reg_7___i169 (.D(write_data_c_8), .SP(clk_c_enable_323), 
            .CK(clk_c), .Q(\key_reg[2] [8]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i169.GSR = "ENABLED";
    FD1P3AX key_reg_7___i170 (.D(write_data_c_9), .SP(clk_c_enable_323), 
            .CK(clk_c), .Q(\key_reg[2] [9]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i170.GSR = "ENABLED";
    FD1P3AX key_reg_7___i171 (.D(write_data_c_10), .SP(clk_c_enable_323), 
            .CK(clk_c), .Q(\key_reg[2] [10]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i171.GSR = "ENABLED";
    FD1P3AX key_reg_7___i172 (.D(write_data_c_11), .SP(clk_c_enable_323), 
            .CK(clk_c), .Q(\key_reg[2] [11]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i172.GSR = "ENABLED";
    FD1P3AX key_reg_7___i173 (.D(write_data_c_12), .SP(clk_c_enable_323), 
            .CK(clk_c), .Q(\key_reg[2] [12]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i173.GSR = "ENABLED";
    FD1P3AX key_reg_7___i174 (.D(write_data_c_13), .SP(clk_c_enable_323), 
            .CK(clk_c), .Q(\key_reg[2] [13]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i174.GSR = "ENABLED";
    FD1P3AX key_reg_7___i175 (.D(write_data_c_14), .SP(clk_c_enable_323), 
            .CK(clk_c), .Q(\key_reg[2] [14]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i175.GSR = "ENABLED";
    FD1P3AX key_reg_7___i176 (.D(write_data_c_15), .SP(clk_c_enable_323), 
            .CK(clk_c), .Q(\key_reg[2] [15]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i176.GSR = "ENABLED";
    FD1P3AX key_reg_7___i177 (.D(write_data_c_16), .SP(clk_c_enable_323), 
            .CK(clk_c), .Q(\key_reg[2] [16]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i177.GSR = "ENABLED";
    FD1P3AX key_reg_7___i178 (.D(write_data_c_17), .SP(clk_c_enable_323), 
            .CK(clk_c), .Q(\key_reg[2] [17]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i178.GSR = "ENABLED";
    FD1P3AX key_reg_7___i179 (.D(write_data_c_18), .SP(clk_c_enable_323), 
            .CK(clk_c), .Q(\key_reg[2] [18]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i179.GSR = "ENABLED";
    FD1P3AX key_reg_7___i180 (.D(write_data_c_19), .SP(clk_c_enable_323), 
            .CK(clk_c), .Q(\key_reg[2] [19]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i180.GSR = "ENABLED";
    FD1P3AX key_reg_7___i181 (.D(write_data_c_20), .SP(clk_c_enable_323), 
            .CK(clk_c), .Q(\key_reg[2] [20]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i181.GSR = "ENABLED";
    FD1P3AX key_reg_7___i182 (.D(write_data_c_21), .SP(clk_c_enable_323), 
            .CK(clk_c), .Q(\key_reg[2] [21]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i182.GSR = "ENABLED";
    FD1P3AX key_reg_7___i183 (.D(write_data_c_22), .SP(clk_c_enable_323), 
            .CK(clk_c), .Q(\key_reg[2] [22]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i183.GSR = "ENABLED";
    FD1P3AX key_reg_7___i184 (.D(write_data_c_23), .SP(clk_c_enable_323), 
            .CK(clk_c), .Q(\key_reg[2] [23]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i184.GSR = "ENABLED";
    FD1P3AX key_reg_7___i185 (.D(write_data_c_24), .SP(clk_c_enable_323), 
            .CK(clk_c), .Q(\key_reg[2] [24]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i185.GSR = "ENABLED";
    FD1P3AX key_reg_7___i186 (.D(write_data_c_25), .SP(clk_c_enable_323), 
            .CK(clk_c), .Q(\key_reg[2] [25]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i186.GSR = "ENABLED";
    FD1P3AX key_reg_7___i187 (.D(write_data_c_26), .SP(clk_c_enable_323), 
            .CK(clk_c), .Q(\key_reg[2] [26]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i187.GSR = "ENABLED";
    FD1P3AX key_reg_7___i188 (.D(write_data_c_27), .SP(clk_c_enable_323), 
            .CK(clk_c), .Q(\key_reg[2] [27]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i188.GSR = "ENABLED";
    FD1P3AX key_reg_7___i189 (.D(write_data_c_28), .SP(clk_c_enable_323), 
            .CK(clk_c), .Q(\key_reg[2] [28]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i189.GSR = "ENABLED";
    FD1P3AX key_reg_7___i190 (.D(write_data_c_29), .SP(clk_c_enable_323), 
            .CK(clk_c), .Q(\key_reg[2] [29]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i190.GSR = "ENABLED";
    FD1P3AX key_reg_7___i191 (.D(write_data_c_30), .SP(clk_c_enable_323), 
            .CK(clk_c), .Q(\key_reg[2] [30]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i191.GSR = "ENABLED";
    FD1P3AX key_reg_7___i192 (.D(write_data_c_31), .SP(clk_c_enable_323), 
            .CK(clk_c), .Q(\key_reg[2] [31]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i192.GSR = "ENABLED";
    FD1P3AX key_reg_7___i193 (.D(write_data_c_0), .SP(clk_c_enable_355), 
            .CK(clk_c), .Q(\key_reg[1] [0]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i193.GSR = "ENABLED";
    FD1P3AX key_reg_7___i194 (.D(write_data_c_1), .SP(clk_c_enable_355), 
            .CK(clk_c), .Q(\key_reg[1] [1]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i194.GSR = "ENABLED";
    FD1P3AX key_reg_7___i195 (.D(write_data_c_2), .SP(clk_c_enable_355), 
            .CK(clk_c), .Q(\key_reg[1] [2]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i195.GSR = "ENABLED";
    FD1P3AX key_reg_7___i196 (.D(write_data_c_3), .SP(clk_c_enable_355), 
            .CK(clk_c), .Q(\key_reg[1] [3]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i196.GSR = "ENABLED";
    FD1P3AX key_reg_7___i197 (.D(write_data_c_4), .SP(clk_c_enable_355), 
            .CK(clk_c), .Q(\key_reg[1] [4]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i197.GSR = "ENABLED";
    FD1P3AX key_reg_7___i198 (.D(write_data_c_5), .SP(clk_c_enable_355), 
            .CK(clk_c), .Q(\key_reg[1] [5]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i198.GSR = "ENABLED";
    FD1P3AX key_reg_7___i199 (.D(write_data_c_6), .SP(clk_c_enable_355), 
            .CK(clk_c), .Q(\key_reg[1] [6]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i199.GSR = "ENABLED";
    FD1P3AX key_reg_7___i200 (.D(write_data_c_7), .SP(clk_c_enable_355), 
            .CK(clk_c), .Q(\key_reg[1] [7]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i200.GSR = "ENABLED";
    FD1P3AX key_reg_7___i201 (.D(write_data_c_8), .SP(clk_c_enable_355), 
            .CK(clk_c), .Q(\key_reg[1] [8]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i201.GSR = "ENABLED";
    FD1P3AX key_reg_7___i202 (.D(write_data_c_9), .SP(clk_c_enable_355), 
            .CK(clk_c), .Q(\key_reg[1] [9]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i202.GSR = "ENABLED";
    FD1P3AX key_reg_7___i203 (.D(write_data_c_10), .SP(clk_c_enable_355), 
            .CK(clk_c), .Q(\key_reg[1] [10]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i203.GSR = "ENABLED";
    FD1P3AX key_reg_7___i204 (.D(write_data_c_11), .SP(clk_c_enable_355), 
            .CK(clk_c), .Q(\key_reg[1] [11]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i204.GSR = "ENABLED";
    FD1P3AX key_reg_7___i205 (.D(write_data_c_12), .SP(clk_c_enable_355), 
            .CK(clk_c), .Q(\key_reg[1] [12]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i205.GSR = "ENABLED";
    FD1P3AX key_reg_7___i206 (.D(write_data_c_13), .SP(clk_c_enable_355), 
            .CK(clk_c), .Q(\key_reg[1] [13]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i206.GSR = "ENABLED";
    FD1P3AX key_reg_7___i207 (.D(write_data_c_14), .SP(clk_c_enable_355), 
            .CK(clk_c), .Q(\key_reg[1] [14]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i207.GSR = "ENABLED";
    FD1P3AX key_reg_7___i208 (.D(write_data_c_15), .SP(clk_c_enable_355), 
            .CK(clk_c), .Q(\key_reg[1] [15]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i208.GSR = "ENABLED";
    FD1P3AX key_reg_7___i209 (.D(write_data_c_16), .SP(clk_c_enable_355), 
            .CK(clk_c), .Q(\key_reg[1] [16]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i209.GSR = "ENABLED";
    FD1P3AX key_reg_7___i210 (.D(write_data_c_17), .SP(clk_c_enable_355), 
            .CK(clk_c), .Q(\key_reg[1] [17]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i210.GSR = "ENABLED";
    FD1P3AX key_reg_7___i211 (.D(write_data_c_18), .SP(clk_c_enable_355), 
            .CK(clk_c), .Q(\key_reg[1] [18]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i211.GSR = "ENABLED";
    FD1P3AX key_reg_7___i212 (.D(write_data_c_19), .SP(clk_c_enable_355), 
            .CK(clk_c), .Q(\key_reg[1] [19]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i212.GSR = "ENABLED";
    FD1P3AX key_reg_7___i213 (.D(write_data_c_20), .SP(clk_c_enable_355), 
            .CK(clk_c), .Q(\key_reg[1] [20]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i213.GSR = "ENABLED";
    FD1P3AX key_reg_7___i214 (.D(write_data_c_21), .SP(clk_c_enable_355), 
            .CK(clk_c), .Q(\key_reg[1] [21]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i214.GSR = "ENABLED";
    FD1P3AX key_reg_7___i215 (.D(write_data_c_22), .SP(clk_c_enable_355), 
            .CK(clk_c), .Q(\key_reg[1] [22]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i215.GSR = "ENABLED";
    FD1P3AX key_reg_7___i216 (.D(write_data_c_23), .SP(clk_c_enable_355), 
            .CK(clk_c), .Q(\key_reg[1] [23]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i216.GSR = "ENABLED";
    FD1P3AX key_reg_7___i217 (.D(write_data_c_24), .SP(clk_c_enable_355), 
            .CK(clk_c), .Q(\key_reg[1] [24]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i217.GSR = "ENABLED";
    FD1P3AX key_reg_7___i218 (.D(write_data_c_25), .SP(clk_c_enable_355), 
            .CK(clk_c), .Q(\key_reg[1] [25]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i218.GSR = "ENABLED";
    FD1P3AX key_reg_7___i219 (.D(write_data_c_26), .SP(clk_c_enable_355), 
            .CK(clk_c), .Q(\key_reg[1] [26]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i219.GSR = "ENABLED";
    FD1P3AX key_reg_7___i220 (.D(write_data_c_27), .SP(clk_c_enable_355), 
            .CK(clk_c), .Q(\key_reg[1] [27]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i220.GSR = "ENABLED";
    FD1P3AX key_reg_7___i221 (.D(write_data_c_28), .SP(clk_c_enable_355), 
            .CK(clk_c), .Q(\key_reg[1] [28]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i221.GSR = "ENABLED";
    FD1P3AX key_reg_7___i222 (.D(write_data_c_29), .SP(clk_c_enable_355), 
            .CK(clk_c), .Q(\key_reg[1] [29]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i222.GSR = "ENABLED";
    FD1P3AX key_reg_7___i223 (.D(write_data_c_30), .SP(clk_c_enable_355), 
            .CK(clk_c), .Q(\key_reg[1] [30]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i223.GSR = "ENABLED";
    FD1P3AX key_reg_7___i224 (.D(write_data_c_31), .SP(clk_c_enable_355), 
            .CK(clk_c), .Q(\key_reg[1] [31]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i224.GSR = "ENABLED";
    FD1P3AX key_reg_7___i225 (.D(write_data_c_0), .SP(clk_c_enable_387), 
            .CK(clk_c), .Q(\key_reg[0] [0]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i225.GSR = "ENABLED";
    FD1P3AX key_reg_7___i226 (.D(write_data_c_1), .SP(clk_c_enable_387), 
            .CK(clk_c), .Q(\key_reg[0] [1]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i226.GSR = "ENABLED";
    FD1P3AX key_reg_7___i227 (.D(write_data_c_2), .SP(clk_c_enable_387), 
            .CK(clk_c), .Q(\key_reg[0] [2]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i227.GSR = "ENABLED";
    FD1P3AX key_reg_7___i228 (.D(write_data_c_3), .SP(clk_c_enable_387), 
            .CK(clk_c), .Q(\key_reg[0] [3]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i228.GSR = "ENABLED";
    FD1P3AX key_reg_7___i229 (.D(write_data_c_4), .SP(clk_c_enable_387), 
            .CK(clk_c), .Q(\key_reg[0] [4]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i229.GSR = "ENABLED";
    FD1P3AX key_reg_7___i230 (.D(write_data_c_5), .SP(clk_c_enable_387), 
            .CK(clk_c), .Q(\key_reg[0] [5]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i230.GSR = "ENABLED";
    FD1P3AX key_reg_7___i231 (.D(write_data_c_6), .SP(clk_c_enable_387), 
            .CK(clk_c), .Q(\key_reg[0] [6]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i231.GSR = "ENABLED";
    FD1P3AX key_reg_7___i232 (.D(write_data_c_7), .SP(clk_c_enable_387), 
            .CK(clk_c), .Q(\key_reg[0] [7]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i232.GSR = "ENABLED";
    FD1P3AX key_reg_7___i233 (.D(write_data_c_8), .SP(clk_c_enable_387), 
            .CK(clk_c), .Q(\key_reg[0] [8]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i233.GSR = "ENABLED";
    FD1P3AX key_reg_7___i234 (.D(write_data_c_9), .SP(clk_c_enable_387), 
            .CK(clk_c), .Q(\key_reg[0] [9]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i234.GSR = "ENABLED";
    FD1P3AX key_reg_7___i235 (.D(write_data_c_10), .SP(clk_c_enable_387), 
            .CK(clk_c), .Q(\key_reg[0] [10]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i235.GSR = "ENABLED";
    FD1P3AX key_reg_7___i236 (.D(write_data_c_11), .SP(clk_c_enable_387), 
            .CK(clk_c), .Q(\key_reg[0] [11]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i236.GSR = "ENABLED";
    FD1P3AX key_reg_7___i237 (.D(write_data_c_12), .SP(clk_c_enable_387), 
            .CK(clk_c), .Q(\key_reg[0] [12]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i237.GSR = "ENABLED";
    FD1P3AX key_reg_7___i238 (.D(write_data_c_13), .SP(clk_c_enable_387), 
            .CK(clk_c), .Q(\key_reg[0] [13]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i238.GSR = "ENABLED";
    FD1P3AX key_reg_7___i239 (.D(write_data_c_14), .SP(clk_c_enable_387), 
            .CK(clk_c), .Q(\key_reg[0] [14]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i239.GSR = "ENABLED";
    FD1P3AX key_reg_7___i240 (.D(write_data_c_15), .SP(clk_c_enable_387), 
            .CK(clk_c), .Q(\key_reg[0] [15]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i240.GSR = "ENABLED";
    FD1P3AX key_reg_7___i241 (.D(write_data_c_16), .SP(clk_c_enable_387), 
            .CK(clk_c), .Q(\key_reg[0] [16]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i241.GSR = "ENABLED";
    FD1P3AX key_reg_7___i242 (.D(write_data_c_17), .SP(clk_c_enable_387), 
            .CK(clk_c), .Q(\key_reg[0] [17]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i242.GSR = "ENABLED";
    FD1P3AX key_reg_7___i243 (.D(write_data_c_18), .SP(clk_c_enable_387), 
            .CK(clk_c), .Q(\key_reg[0] [18]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i243.GSR = "ENABLED";
    FD1P3AX key_reg_7___i244 (.D(write_data_c_19), .SP(clk_c_enable_387), 
            .CK(clk_c), .Q(\key_reg[0] [19]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i244.GSR = "ENABLED";
    FD1P3AX key_reg_7___i245 (.D(write_data_c_20), .SP(clk_c_enable_387), 
            .CK(clk_c), .Q(\key_reg[0] [20]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i245.GSR = "ENABLED";
    FD1P3AX key_reg_7___i246 (.D(write_data_c_21), .SP(clk_c_enable_387), 
            .CK(clk_c), .Q(\key_reg[0] [21]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i246.GSR = "ENABLED";
    FD1P3AX key_reg_7___i247 (.D(write_data_c_22), .SP(clk_c_enable_387), 
            .CK(clk_c), .Q(\key_reg[0] [22]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i247.GSR = "ENABLED";
    FD1P3AX key_reg_7___i248 (.D(write_data_c_23), .SP(clk_c_enable_387), 
            .CK(clk_c), .Q(\key_reg[0] [23]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i248.GSR = "ENABLED";
    FD1P3AX key_reg_7___i249 (.D(write_data_c_24), .SP(clk_c_enable_387), 
            .CK(clk_c), .Q(\key_reg[0] [24]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i249.GSR = "ENABLED";
    FD1P3AX key_reg_7___i250 (.D(write_data_c_25), .SP(clk_c_enable_387), 
            .CK(clk_c), .Q(\key_reg[0] [25]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i250.GSR = "ENABLED";
    FD1P3AX key_reg_7___i251 (.D(write_data_c_26), .SP(clk_c_enable_387), 
            .CK(clk_c), .Q(\key_reg[0] [26]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i251.GSR = "ENABLED";
    FD1P3AX key_reg_7___i252 (.D(write_data_c_27), .SP(clk_c_enable_387), 
            .CK(clk_c), .Q(\key_reg[0] [27]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i252.GSR = "ENABLED";
    FD1P3AX key_reg_7___i253 (.D(write_data_c_28), .SP(clk_c_enable_387), 
            .CK(clk_c), .Q(\key_reg[0] [28]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i253.GSR = "ENABLED";
    FD1P3AX key_reg_7___i254 (.D(write_data_c_29), .SP(clk_c_enable_387), 
            .CK(clk_c), .Q(\key_reg[0] [29]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i254.GSR = "ENABLED";
    FD1P3AX key_reg_7___i255 (.D(write_data_c_30), .SP(clk_c_enable_387), 
            .CK(clk_c), .Q(\key_reg[0] [30]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i255.GSR = "ENABLED";
    FD1P3AX key_reg_7___i256 (.D(write_data_c_31), .SP(clk_c_enable_387), 
            .CK(clk_c), .Q(\key_reg[0] [31]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam key_reg_7___i256.GSR = "ENABLED";
    LUT4 i25785_then_3_lut (.A(result_reg[72]), .B(address_c_1), .C(result_reg[8]), 
         .Z(n33996)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i25785_then_3_lut.init = 16'he2e2;
    LUT4 i27886_2_lut_4_lut_4_lut (.A(n33949), .B(n33857), .C(n28824), 
         .D(n33910), .Z(clk_c_enable_2540)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i27886_2_lut_4_lut_4_lut.init = 16'h0040;
    LUT4 i27855_2_lut_4_lut_4_lut (.A(n33940), .B(n33857), .C(n28824), 
         .D(n33910), .Z(clk_c_enable_2508)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i27855_2_lut_4_lut_4_lut.init = 16'h0040;
    LUT4 i27884_2_lut_4_lut_4_lut (.A(n33946), .B(n33857), .C(n28824), 
         .D(n33910), .Z(clk_c_enable_2476)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i27884_2_lut_4_lut_4_lut.init = 16'h0040;
    LUT4 i25785_else_3_lut (.A(result_reg[104]), .B(address_c_1), .C(result_reg[40]), 
         .Z(n33995)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i25785_else_3_lut.init = 16'he2e2;
    LUT4 i25788_then_3_lut (.A(result_reg[73]), .B(address_c_1), .C(result_reg[9]), 
         .Z(n33999)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i25788_then_3_lut.init = 16'he2e2;
    LUT4 i25788_else_3_lut (.A(result_reg[105]), .B(address_c_1), .C(result_reg[41]), 
         .Z(n33998)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i25788_else_3_lut.init = 16'he2e2;
    PFUMX i29048 (.BLUT(n33998), .ALUT(n33999), .C0(address_c_0), .Z(n34000));
    LUT4 i25791_then_3_lut (.A(result_reg[74]), .B(address_c_1), .C(result_reg[10]), 
         .Z(n34002)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i25791_then_3_lut.init = 16'he2e2;
    LUT4 i25791_else_3_lut (.A(result_reg[106]), .B(address_c_1), .C(result_reg[42]), 
         .Z(n34001)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i25791_else_3_lut.init = 16'he2e2;
    PFUMX i29046 (.BLUT(n33995), .ALUT(n33996), .C0(address_c_0), .Z(n33997));
    LUT4 i15188_3_lut (.A(key_mem_ctrl_new_2__N_4928[0]), .B(aes_core_ctrl_reg[1]), 
         .C(aes_core_ctrl_reg[0]), .Z(init_state)) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(274[7] 331[14])
    defparam i15188_3_lut.init = 16'h3232;
    FD1P3AX block_reg_3___i2 (.D(write_data_c_1), .SP(clk_c_enable_2444), 
            .CK(clk_c), .Q(\block_reg[3] [1]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i2.GSR = "ENABLED";
    FD1P3AX block_reg_3___i3 (.D(write_data_c_2), .SP(clk_c_enable_2444), 
            .CK(clk_c), .Q(\block_reg[3] [2]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i3.GSR = "ENABLED";
    FD1P3AX block_reg_3___i4 (.D(write_data_c_3), .SP(clk_c_enable_2444), 
            .CK(clk_c), .Q(\block_reg[3] [3]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i4.GSR = "ENABLED";
    FD1P3AX block_reg_3___i5 (.D(write_data_c_4), .SP(clk_c_enable_2444), 
            .CK(clk_c), .Q(\block_reg[3] [4]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i5.GSR = "ENABLED";
    FD1P3AX block_reg_3___i6 (.D(write_data_c_5), .SP(clk_c_enable_2444), 
            .CK(clk_c), .Q(\block_reg[3] [5]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i6.GSR = "ENABLED";
    FD1P3AX block_reg_3___i7 (.D(write_data_c_6), .SP(clk_c_enable_2444), 
            .CK(clk_c), .Q(\block_reg[3] [6]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i7.GSR = "ENABLED";
    FD1P3AX block_reg_3___i8 (.D(write_data_c_7), .SP(clk_c_enable_2444), 
            .CK(clk_c), .Q(\block_reg[3] [7]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i8.GSR = "ENABLED";
    FD1P3AX block_reg_3___i9 (.D(write_data_c_8), .SP(clk_c_enable_2444), 
            .CK(clk_c), .Q(\block_reg[3] [8]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i9.GSR = "ENABLED";
    FD1P3AX block_reg_3___i10 (.D(write_data_c_9), .SP(clk_c_enable_2444), 
            .CK(clk_c), .Q(\block_reg[3] [9]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i10.GSR = "ENABLED";
    FD1P3AX block_reg_3___i11 (.D(write_data_c_10), .SP(clk_c_enable_2444), 
            .CK(clk_c), .Q(\block_reg[3] [10]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i11.GSR = "ENABLED";
    FD1P3AX block_reg_3___i12 (.D(write_data_c_11), .SP(clk_c_enable_2444), 
            .CK(clk_c), .Q(\block_reg[3] [11]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i12.GSR = "ENABLED";
    FD1P3AX block_reg_3___i13 (.D(write_data_c_12), .SP(clk_c_enable_2444), 
            .CK(clk_c), .Q(\block_reg[3] [12]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i13.GSR = "ENABLED";
    FD1P3AX block_reg_3___i14 (.D(write_data_c_13), .SP(clk_c_enable_2444), 
            .CK(clk_c), .Q(\block_reg[3] [13]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i14.GSR = "ENABLED";
    FD1P3AX block_reg_3___i15 (.D(write_data_c_14), .SP(clk_c_enable_2444), 
            .CK(clk_c), .Q(\block_reg[3] [14]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i15.GSR = "ENABLED";
    FD1P3AX block_reg_3___i16 (.D(write_data_c_15), .SP(clk_c_enable_2444), 
            .CK(clk_c), .Q(\block_reg[3] [15]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i16.GSR = "ENABLED";
    FD1P3AX block_reg_3___i17 (.D(write_data_c_16), .SP(clk_c_enable_2444), 
            .CK(clk_c), .Q(\block_reg[3] [16]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i17.GSR = "ENABLED";
    FD1P3AX block_reg_3___i18 (.D(write_data_c_17), .SP(clk_c_enable_2444), 
            .CK(clk_c), .Q(\block_reg[3] [17]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i18.GSR = "ENABLED";
    FD1P3AX block_reg_3___i19 (.D(write_data_c_18), .SP(clk_c_enable_2444), 
            .CK(clk_c), .Q(\block_reg[3] [18]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i19.GSR = "ENABLED";
    FD1P3AX block_reg_3___i20 (.D(write_data_c_19), .SP(clk_c_enable_2444), 
            .CK(clk_c), .Q(\block_reg[3] [19]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i20.GSR = "ENABLED";
    FD1P3AX block_reg_3___i21 (.D(write_data_c_20), .SP(clk_c_enable_2444), 
            .CK(clk_c), .Q(\block_reg[3] [20]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i21.GSR = "ENABLED";
    FD1P3AX block_reg_3___i22 (.D(write_data_c_21), .SP(clk_c_enable_2444), 
            .CK(clk_c), .Q(\block_reg[3] [21]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i22.GSR = "ENABLED";
    FD1P3AX block_reg_3___i23 (.D(write_data_c_22), .SP(clk_c_enable_2444), 
            .CK(clk_c), .Q(\block_reg[3] [22]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i23.GSR = "ENABLED";
    FD1P3AX block_reg_3___i24 (.D(write_data_c_23), .SP(clk_c_enable_2444), 
            .CK(clk_c), .Q(\block_reg[3] [23]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i24.GSR = "ENABLED";
    FD1P3AX block_reg_3___i25 (.D(write_data_c_24), .SP(clk_c_enable_2444), 
            .CK(clk_c), .Q(\block_reg[3] [24]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i25.GSR = "ENABLED";
    FD1P3AX block_reg_3___i26 (.D(write_data_c_25), .SP(clk_c_enable_2444), 
            .CK(clk_c), .Q(\block_reg[3] [25]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i26.GSR = "ENABLED";
    FD1P3AX block_reg_3___i27 (.D(write_data_c_26), .SP(clk_c_enable_2444), 
            .CK(clk_c), .Q(\block_reg[3] [26]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i27.GSR = "ENABLED";
    FD1P3AX block_reg_3___i28 (.D(write_data_c_27), .SP(clk_c_enable_2444), 
            .CK(clk_c), .Q(\block_reg[3] [27]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i28.GSR = "ENABLED";
    FD1P3AX block_reg_3___i29 (.D(write_data_c_28), .SP(clk_c_enable_2444), 
            .CK(clk_c), .Q(\block_reg[3] [28]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i29.GSR = "ENABLED";
    FD1P3AX block_reg_3___i30 (.D(write_data_c_29), .SP(clk_c_enable_2444), 
            .CK(clk_c), .Q(\block_reg[3] [29]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i30.GSR = "ENABLED";
    FD1P3AX block_reg_3___i31 (.D(write_data_c_30), .SP(clk_c_enable_2444), 
            .CK(clk_c), .Q(\block_reg[3] [30]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i31.GSR = "ENABLED";
    FD1P3AX block_reg_3___i32 (.D(write_data_c_31), .SP(clk_c_enable_2444), 
            .CK(clk_c), .Q(\block_reg[3] [31]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i32.GSR = "ENABLED";
    FD1P3AX block_reg_3___i33 (.D(write_data_c_0), .SP(clk_c_enable_2476), 
            .CK(clk_c), .Q(\block_reg[2] [0]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i33.GSR = "ENABLED";
    FD1P3AX block_reg_3___i34 (.D(write_data_c_1), .SP(clk_c_enable_2476), 
            .CK(clk_c), .Q(\block_reg[2] [1]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i34.GSR = "ENABLED";
    FD1P3AX block_reg_3___i35 (.D(write_data_c_2), .SP(clk_c_enable_2476), 
            .CK(clk_c), .Q(\block_reg[2] [2]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i35.GSR = "ENABLED";
    FD1P3AX block_reg_3___i36 (.D(write_data_c_3), .SP(clk_c_enable_2476), 
            .CK(clk_c), .Q(\block_reg[2] [3]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i36.GSR = "ENABLED";
    FD1P3AX block_reg_3___i37 (.D(write_data_c_4), .SP(clk_c_enable_2476), 
            .CK(clk_c), .Q(\block_reg[2] [4]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i37.GSR = "ENABLED";
    FD1P3AX block_reg_3___i38 (.D(write_data_c_5), .SP(clk_c_enable_2476), 
            .CK(clk_c), .Q(\block_reg[2] [5]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i38.GSR = "ENABLED";
    FD1P3AX block_reg_3___i39 (.D(write_data_c_6), .SP(clk_c_enable_2476), 
            .CK(clk_c), .Q(\block_reg[2] [6]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i39.GSR = "ENABLED";
    FD1P3AX block_reg_3___i40 (.D(write_data_c_7), .SP(clk_c_enable_2476), 
            .CK(clk_c), .Q(\block_reg[2] [7]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i40.GSR = "ENABLED";
    FD1P3AX block_reg_3___i41 (.D(write_data_c_8), .SP(clk_c_enable_2476), 
            .CK(clk_c), .Q(\block_reg[2] [8]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i41.GSR = "ENABLED";
    FD1P3AX block_reg_3___i42 (.D(write_data_c_9), .SP(clk_c_enable_2476), 
            .CK(clk_c), .Q(\block_reg[2] [9]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i42.GSR = "ENABLED";
    FD1P3AX block_reg_3___i43 (.D(write_data_c_10), .SP(clk_c_enable_2476), 
            .CK(clk_c), .Q(\block_reg[2] [10]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i43.GSR = "ENABLED";
    FD1P3AX block_reg_3___i44 (.D(write_data_c_11), .SP(clk_c_enable_2476), 
            .CK(clk_c), .Q(\block_reg[2] [11]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i44.GSR = "ENABLED";
    FD1P3AX block_reg_3___i45 (.D(write_data_c_12), .SP(clk_c_enable_2476), 
            .CK(clk_c), .Q(\block_reg[2] [12]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i45.GSR = "ENABLED";
    FD1P3AX block_reg_3___i46 (.D(write_data_c_13), .SP(clk_c_enable_2476), 
            .CK(clk_c), .Q(\block_reg[2] [13]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i46.GSR = "ENABLED";
    FD1P3AX block_reg_3___i47 (.D(write_data_c_14), .SP(clk_c_enable_2476), 
            .CK(clk_c), .Q(\block_reg[2] [14]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i47.GSR = "ENABLED";
    FD1P3AX block_reg_3___i48 (.D(write_data_c_15), .SP(clk_c_enable_2476), 
            .CK(clk_c), .Q(\block_reg[2] [15]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i48.GSR = "ENABLED";
    FD1P3AX block_reg_3___i49 (.D(write_data_c_16), .SP(clk_c_enable_2476), 
            .CK(clk_c), .Q(\block_reg[2] [16]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i49.GSR = "ENABLED";
    FD1P3AX block_reg_3___i50 (.D(write_data_c_17), .SP(clk_c_enable_2476), 
            .CK(clk_c), .Q(\block_reg[2] [17]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i50.GSR = "ENABLED";
    FD1P3AX block_reg_3___i51 (.D(write_data_c_18), .SP(clk_c_enable_2476), 
            .CK(clk_c), .Q(\block_reg[2] [18]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i51.GSR = "ENABLED";
    FD1P3AX block_reg_3___i52 (.D(write_data_c_19), .SP(clk_c_enable_2476), 
            .CK(clk_c), .Q(\block_reg[2] [19]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i52.GSR = "ENABLED";
    FD1P3AX block_reg_3___i53 (.D(write_data_c_20), .SP(clk_c_enable_2476), 
            .CK(clk_c), .Q(\block_reg[2] [20]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i53.GSR = "ENABLED";
    FD1P3AX block_reg_3___i54 (.D(write_data_c_21), .SP(clk_c_enable_2476), 
            .CK(clk_c), .Q(\block_reg[2] [21]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i54.GSR = "ENABLED";
    FD1P3AX block_reg_3___i55 (.D(write_data_c_22), .SP(clk_c_enable_2476), 
            .CK(clk_c), .Q(\block_reg[2] [22]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i55.GSR = "ENABLED";
    FD1P3AX block_reg_3___i56 (.D(write_data_c_23), .SP(clk_c_enable_2476), 
            .CK(clk_c), .Q(\block_reg[2] [23]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i56.GSR = "ENABLED";
    FD1P3AX block_reg_3___i57 (.D(write_data_c_24), .SP(clk_c_enable_2476), 
            .CK(clk_c), .Q(\block_reg[2] [24]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i57.GSR = "ENABLED";
    FD1P3AX block_reg_3___i58 (.D(write_data_c_25), .SP(clk_c_enable_2476), 
            .CK(clk_c), .Q(\block_reg[2] [25]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i58.GSR = "ENABLED";
    FD1P3AX block_reg_3___i59 (.D(write_data_c_26), .SP(clk_c_enable_2476), 
            .CK(clk_c), .Q(\block_reg[2] [26]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i59.GSR = "ENABLED";
    FD1P3AX block_reg_3___i60 (.D(write_data_c_27), .SP(clk_c_enable_2476), 
            .CK(clk_c), .Q(\block_reg[2] [27]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i60.GSR = "ENABLED";
    FD1P3AX block_reg_3___i61 (.D(write_data_c_28), .SP(clk_c_enable_2476), 
            .CK(clk_c), .Q(\block_reg[2] [28]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i61.GSR = "ENABLED";
    FD1P3AX block_reg_3___i62 (.D(write_data_c_29), .SP(clk_c_enable_2476), 
            .CK(clk_c), .Q(\block_reg[2] [29]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i62.GSR = "ENABLED";
    FD1P3AX block_reg_3___i63 (.D(write_data_c_30), .SP(clk_c_enable_2476), 
            .CK(clk_c), .Q(\block_reg[2] [30]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i63.GSR = "ENABLED";
    FD1P3AX block_reg_3___i64 (.D(write_data_c_31), .SP(clk_c_enable_2476), 
            .CK(clk_c), .Q(\block_reg[2] [31]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i64.GSR = "ENABLED";
    FD1P3AX block_reg_3___i65 (.D(write_data_c_0), .SP(clk_c_enable_2508), 
            .CK(clk_c), .Q(\block_reg[1] [0]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i65.GSR = "ENABLED";
    FD1P3AX block_reg_3___i66 (.D(write_data_c_1), .SP(clk_c_enable_2508), 
            .CK(clk_c), .Q(\block_reg[1] [1]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i66.GSR = "ENABLED";
    FD1P3AX block_reg_3___i67 (.D(write_data_c_2), .SP(clk_c_enable_2508), 
            .CK(clk_c), .Q(\block_reg[1] [2]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i67.GSR = "ENABLED";
    FD1P3AX block_reg_3___i68 (.D(write_data_c_3), .SP(clk_c_enable_2508), 
            .CK(clk_c), .Q(\block_reg[1] [3]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i68.GSR = "ENABLED";
    FD1P3AX block_reg_3___i69 (.D(write_data_c_4), .SP(clk_c_enable_2508), 
            .CK(clk_c), .Q(\block_reg[1] [4]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i69.GSR = "ENABLED";
    FD1P3AX block_reg_3___i70 (.D(write_data_c_5), .SP(clk_c_enable_2508), 
            .CK(clk_c), .Q(\block_reg[1] [5]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i70.GSR = "ENABLED";
    FD1P3AX block_reg_3___i71 (.D(write_data_c_6), .SP(clk_c_enable_2508), 
            .CK(clk_c), .Q(\block_reg[1] [6]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i71.GSR = "ENABLED";
    FD1P3AX block_reg_3___i72 (.D(write_data_c_7), .SP(clk_c_enable_2508), 
            .CK(clk_c), .Q(\block_reg[1] [7]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i72.GSR = "ENABLED";
    FD1P3AX block_reg_3___i73 (.D(write_data_c_8), .SP(clk_c_enable_2508), 
            .CK(clk_c), .Q(\block_reg[1] [8]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i73.GSR = "ENABLED";
    FD1P3AX block_reg_3___i74 (.D(write_data_c_9), .SP(clk_c_enable_2508), 
            .CK(clk_c), .Q(\block_reg[1] [9]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i74.GSR = "ENABLED";
    FD1P3AX block_reg_3___i75 (.D(write_data_c_10), .SP(clk_c_enable_2508), 
            .CK(clk_c), .Q(\block_reg[1] [10]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i75.GSR = "ENABLED";
    FD1P3AX block_reg_3___i76 (.D(write_data_c_11), .SP(clk_c_enable_2508), 
            .CK(clk_c), .Q(\block_reg[1] [11]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i76.GSR = "ENABLED";
    FD1P3AX block_reg_3___i77 (.D(write_data_c_12), .SP(clk_c_enable_2508), 
            .CK(clk_c), .Q(\block_reg[1] [12]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i77.GSR = "ENABLED";
    FD1P3AX block_reg_3___i78 (.D(write_data_c_13), .SP(clk_c_enable_2508), 
            .CK(clk_c), .Q(\block_reg[1] [13]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i78.GSR = "ENABLED";
    FD1P3AX block_reg_3___i79 (.D(write_data_c_14), .SP(clk_c_enable_2508), 
            .CK(clk_c), .Q(\block_reg[1] [14]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i79.GSR = "ENABLED";
    FD1P3AX block_reg_3___i80 (.D(write_data_c_15), .SP(clk_c_enable_2508), 
            .CK(clk_c), .Q(\block_reg[1] [15]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i80.GSR = "ENABLED";
    FD1P3AX block_reg_3___i81 (.D(write_data_c_16), .SP(clk_c_enable_2508), 
            .CK(clk_c), .Q(\block_reg[1] [16]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i81.GSR = "ENABLED";
    FD1P3AX block_reg_3___i82 (.D(write_data_c_17), .SP(clk_c_enable_2508), 
            .CK(clk_c), .Q(\block_reg[1] [17]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i82.GSR = "ENABLED";
    FD1P3AX block_reg_3___i83 (.D(write_data_c_18), .SP(clk_c_enable_2508), 
            .CK(clk_c), .Q(\block_reg[1] [18]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i83.GSR = "ENABLED";
    FD1P3AX block_reg_3___i84 (.D(write_data_c_19), .SP(clk_c_enable_2508), 
            .CK(clk_c), .Q(\block_reg[1] [19]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i84.GSR = "ENABLED";
    FD1P3AX block_reg_3___i85 (.D(write_data_c_20), .SP(clk_c_enable_2508), 
            .CK(clk_c), .Q(\block_reg[1] [20]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i85.GSR = "ENABLED";
    FD1P3AX block_reg_3___i86 (.D(write_data_c_21), .SP(clk_c_enable_2508), 
            .CK(clk_c), .Q(\block_reg[1] [21]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i86.GSR = "ENABLED";
    FD1P3AX block_reg_3___i87 (.D(write_data_c_22), .SP(clk_c_enable_2508), 
            .CK(clk_c), .Q(\block_reg[1] [22]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i87.GSR = "ENABLED";
    FD1P3AX block_reg_3___i88 (.D(write_data_c_23), .SP(clk_c_enable_2508), 
            .CK(clk_c), .Q(\block_reg[1] [23]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i88.GSR = "ENABLED";
    FD1P3AX block_reg_3___i89 (.D(write_data_c_24), .SP(clk_c_enable_2508), 
            .CK(clk_c), .Q(\block_reg[1] [24]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i89.GSR = "ENABLED";
    FD1P3AX block_reg_3___i90 (.D(write_data_c_25), .SP(clk_c_enable_2508), 
            .CK(clk_c), .Q(\block_reg[1] [25]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i90.GSR = "ENABLED";
    FD1P3AX block_reg_3___i91 (.D(write_data_c_26), .SP(clk_c_enable_2508), 
            .CK(clk_c), .Q(\block_reg[1] [26]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i91.GSR = "ENABLED";
    FD1P3AX block_reg_3___i92 (.D(write_data_c_27), .SP(clk_c_enable_2508), 
            .CK(clk_c), .Q(\block_reg[1] [27]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i92.GSR = "ENABLED";
    FD1P3AX block_reg_3___i93 (.D(write_data_c_28), .SP(clk_c_enable_2508), 
            .CK(clk_c), .Q(\block_reg[1] [28]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i93.GSR = "ENABLED";
    FD1P3AX block_reg_3___i94 (.D(write_data_c_29), .SP(clk_c_enable_2508), 
            .CK(clk_c), .Q(\block_reg[1] [29]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i94.GSR = "ENABLED";
    FD1P3AX block_reg_3___i95 (.D(write_data_c_30), .SP(clk_c_enable_2508), 
            .CK(clk_c), .Q(\block_reg[1] [30]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i95.GSR = "ENABLED";
    FD1P3AX block_reg_3___i96 (.D(write_data_c_31), .SP(clk_c_enable_2508), 
            .CK(clk_c), .Q(\block_reg[1] [31]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i96.GSR = "ENABLED";
    FD1P3AX block_reg_3___i97 (.D(write_data_c_0), .SP(clk_c_enable_2540), 
            .CK(clk_c), .Q(\block_reg[0] [0]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i97.GSR = "ENABLED";
    FD1P3AX block_reg_3___i98 (.D(write_data_c_1), .SP(clk_c_enable_2540), 
            .CK(clk_c), .Q(\block_reg[0] [1]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i98.GSR = "ENABLED";
    FD1P3AX block_reg_3___i99 (.D(write_data_c_2), .SP(clk_c_enable_2540), 
            .CK(clk_c), .Q(\block_reg[0] [2]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i99.GSR = "ENABLED";
    FD1P3AX block_reg_3___i100 (.D(write_data_c_3), .SP(clk_c_enable_2540), 
            .CK(clk_c), .Q(\block_reg[0] [3]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i100.GSR = "ENABLED";
    FD1P3AX block_reg_3___i101 (.D(write_data_c_4), .SP(clk_c_enable_2540), 
            .CK(clk_c), .Q(\block_reg[0] [4]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i101.GSR = "ENABLED";
    FD1P3AX block_reg_3___i102 (.D(write_data_c_5), .SP(clk_c_enable_2540), 
            .CK(clk_c), .Q(\block_reg[0] [5]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i102.GSR = "ENABLED";
    FD1P3AX block_reg_3___i103 (.D(write_data_c_6), .SP(clk_c_enable_2540), 
            .CK(clk_c), .Q(\block_reg[0] [6]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i103.GSR = "ENABLED";
    FD1P3AX block_reg_3___i104 (.D(write_data_c_7), .SP(clk_c_enable_2540), 
            .CK(clk_c), .Q(\block_reg[0] [7]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i104.GSR = "ENABLED";
    FD1P3AX block_reg_3___i105 (.D(write_data_c_8), .SP(clk_c_enable_2540), 
            .CK(clk_c), .Q(\block_reg[0] [8]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i105.GSR = "ENABLED";
    FD1P3AX block_reg_3___i106 (.D(write_data_c_9), .SP(clk_c_enable_2540), 
            .CK(clk_c), .Q(\block_reg[0] [9]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i106.GSR = "ENABLED";
    FD1P3AX block_reg_3___i107 (.D(write_data_c_10), .SP(clk_c_enable_2540), 
            .CK(clk_c), .Q(\block_reg[0] [10]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i107.GSR = "ENABLED";
    FD1P3AX block_reg_3___i108 (.D(write_data_c_11), .SP(clk_c_enable_2540), 
            .CK(clk_c), .Q(\block_reg[0] [11]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i108.GSR = "ENABLED";
    FD1P3AX block_reg_3___i109 (.D(write_data_c_12), .SP(clk_c_enable_2540), 
            .CK(clk_c), .Q(\block_reg[0] [12]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i109.GSR = "ENABLED";
    FD1P3AX block_reg_3___i110 (.D(write_data_c_13), .SP(clk_c_enable_2540), 
            .CK(clk_c), .Q(\block_reg[0] [13]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i110.GSR = "ENABLED";
    FD1P3AX block_reg_3___i111 (.D(write_data_c_14), .SP(clk_c_enable_2540), 
            .CK(clk_c), .Q(\block_reg[0] [14]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i111.GSR = "ENABLED";
    FD1P3AX block_reg_3___i112 (.D(write_data_c_15), .SP(clk_c_enable_2540), 
            .CK(clk_c), .Q(\block_reg[0] [15]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i112.GSR = "ENABLED";
    FD1P3AX block_reg_3___i113 (.D(write_data_c_16), .SP(clk_c_enable_2540), 
            .CK(clk_c), .Q(\block_reg[0] [16]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i113.GSR = "ENABLED";
    FD1P3AX block_reg_3___i114 (.D(write_data_c_17), .SP(clk_c_enable_2540), 
            .CK(clk_c), .Q(\block_reg[0] [17]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i114.GSR = "ENABLED";
    FD1P3AX block_reg_3___i115 (.D(write_data_c_18), .SP(clk_c_enable_2540), 
            .CK(clk_c), .Q(\block_reg[0] [18]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i115.GSR = "ENABLED";
    FD1P3AX block_reg_3___i116 (.D(write_data_c_19), .SP(clk_c_enable_2540), 
            .CK(clk_c), .Q(\block_reg[0] [19]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i116.GSR = "ENABLED";
    FD1P3AX block_reg_3___i117 (.D(write_data_c_20), .SP(clk_c_enable_2540), 
            .CK(clk_c), .Q(\block_reg[0] [20]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i117.GSR = "ENABLED";
    FD1P3AX block_reg_3___i118 (.D(write_data_c_21), .SP(clk_c_enable_2540), 
            .CK(clk_c), .Q(\block_reg[0] [21]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i118.GSR = "ENABLED";
    FD1P3AX block_reg_3___i119 (.D(write_data_c_22), .SP(clk_c_enable_2540), 
            .CK(clk_c), .Q(\block_reg[0] [22]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i119.GSR = "ENABLED";
    FD1P3AX block_reg_3___i120 (.D(write_data_c_23), .SP(clk_c_enable_2540), 
            .CK(clk_c), .Q(\block_reg[0] [23]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i120.GSR = "ENABLED";
    FD1P3AX block_reg_3___i121 (.D(write_data_c_24), .SP(clk_c_enable_2540), 
            .CK(clk_c), .Q(\block_reg[0] [24]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i121.GSR = "ENABLED";
    FD1P3AX block_reg_3___i122 (.D(write_data_c_25), .SP(clk_c_enable_2540), 
            .CK(clk_c), .Q(\block_reg[0] [25]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i122.GSR = "ENABLED";
    FD1P3AX block_reg_3___i123 (.D(write_data_c_26), .SP(clk_c_enable_2540), 
            .CK(clk_c), .Q(\block_reg[0] [26]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i123.GSR = "ENABLED";
    FD1P3AX block_reg_3___i124 (.D(write_data_c_27), .SP(clk_c_enable_2540), 
            .CK(clk_c), .Q(\block_reg[0] [27]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i124.GSR = "ENABLED";
    FD1P3AX block_reg_3___i125 (.D(write_data_c_28), .SP(clk_c_enable_2540), 
            .CK(clk_c), .Q(\block_reg[0] [28]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i125.GSR = "ENABLED";
    FD1P3AX block_reg_3___i126 (.D(write_data_c_29), .SP(clk_c_enable_2540), 
            .CK(clk_c), .Q(\block_reg[0] [29]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i126.GSR = "ENABLED";
    FD1P3AX block_reg_3___i127 (.D(write_data_c_30), .SP(clk_c_enable_2540), 
            .CK(clk_c), .Q(\block_reg[0] [30]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i127.GSR = "ENABLED";
    FD1P3AX block_reg_3___i128 (.D(write_data_c_31), .SP(clk_c_enable_2540), 
            .CK(clk_c), .Q(\block_reg[0] [31]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam block_reg_3___i128.GSR = "ENABLED";
    PFUMX i29044 (.BLUT(n33992), .ALUT(n33993), .C0(address_c_0), .Z(n33994));
    FD1S3IX next_reg_104 (.D(n10461), .CK(clk_c), .CD(n13203), .Q(aes_core_ctrl_new_1__N_858[1]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam next_reg_104.GSR = "ENABLED";
    FD1S3IX init_reg_103 (.D(n10461), .CK(clk_c), .CD(n13202), .Q(key_mem_ctrl_new_2__N_4928[0]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam init_reg_103.GSR = "ENABLED";
    GSR GSR_INST (.GSR(reset_n_c));
    PFUMX i29042 (.BLUT(n33989), .ALUT(n33990), .C0(address_c_0), .Z(n33991));
    PFUMX i29040 (.BLUT(n33986), .ALUT(n33987), .C0(address_c_0), .Z(n33988));
    PFUMX i29038 (.BLUT(n33983), .ALUT(n33984), .C0(address_c_0), .Z(n33985));
    PFUMX i29036 (.BLUT(n33980), .ALUT(n33981), .C0(address_c_1), .Z(read_data_c_27));
    PFUMX i29034 (.BLUT(n33977), .ALUT(n33978), .C0(address_c_1), .Z(read_data_c_15));
    PFUMX i29032 (.BLUT(n33974), .ALUT(n33975), .C0(address_c_1), .Z(read_data_c_25));
    PFUMX i29030 (.BLUT(n33971), .ALUT(n33972), .C0(address_c_1), .Z(read_data_c_31));
    PFUMX i29028 (.BLUT(n33968), .ALUT(n33969), .C0(address_c_1), .Z(read_data_c_7));
    PFUMX i29026 (.BLUT(n33965), .ALUT(n33966), .C0(address_c_1), .Z(read_data_c_26));
    PFUMX i29024 (.BLUT(n33962), .ALUT(n33963), .C0(address_c_1), .Z(read_data_c_23));
    LUT4 i2_3_lut_rep_546_4_lut (.A(n33939), .B(address_c_3), .C(address_c_4), 
         .D(n15362), .Z(n33850)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i2_3_lut_rep_546_4_lut.init = 16'h0020;
    LUT4 i2_3_lut_4_lut_adj_851 (.A(encdec_reg), .B(n33942), .C(n149), 
         .D(n33909), .Z(dec_ctrl_we)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i2_3_lut_4_lut_adj_851.init = 16'hfff4;
    LUT4 i1_3_lut_4_lut (.A(encdec_reg), .B(n33942), .C(dec_round_nr[0]), 
         .D(n149), .Z(round_ctr_new[0])) /* synthesis lut_function=(!(A (C+!(D))+!A (B+(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut.init = 16'h0b00;
    LUT4 i1_3_lut_4_lut_adj_852 (.A(encdec_reg), .B(n33942), .C(n149), 
         .D(n14939), .Z(round_ctr_new[3])) /* synthesis lut_function=(A (C (D))+!A (B+(C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_adj_852.init = 16'hf444;
    PFUMX i29022 (.BLUT(n33959), .ALUT(n33960), .C0(address_c_1), .Z(read_data_c_6));
    LUT4 mux_194_Mux_0_i3_3_lut_4_lut (.A(n33948), .B(aes_core_ctrl_reg[0]), 
         .C(aes_core_ctrl_reg[1]), .D(n1), .Z(ready_we)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(274[7] 331[14])
    defparam mux_194_Mux_0_i3_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_196_Mux_0_i3_4_lut_4_lut (.A(n33948), .B(aes_core_ctrl_reg[0]), 
         .C(aes_core_ctrl_reg[1]), .D(n33947), .Z(result_valid_we)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A !(B+(C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(274[7] 331[14])
    defparam mux_196_Mux_0_i3_4_lut_4_lut.init = 16'h8380;
    LUT4 i2_2_lut_3_lut (.A(n33948), .B(aes_core_ctrl_reg[0]), .C(aes_core_ctrl_reg[1]), 
         .Z(result_valid_new)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(274[7] 331[14])
    defparam i2_2_lut_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n15362), .B(n33910), .C(address_c_1), 
         .D(address_c_3), .Z(n28830)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(49[33:40])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i1_2_lut_3_lut_4_lut_adj_853 (.A(n15362), .B(n33910), .C(n33949), 
         .D(address_c_3), .Z(n37)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(49[33:40])
    defparam i1_2_lut_3_lut_4_lut_adj_853.init = 16'hfffe;
    LUT4 i2_3_lut_4_lut_adj_854 (.A(n15362), .B(n33910), .C(address_c_3), 
         .D(n33941), .Z(n25954)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(49[33:40])
    defparam i2_3_lut_4_lut_adj_854.init = 16'hfffe;
    LUT4 i15233_2_lut_3_lut_4_lut (.A(n15362), .B(n33910), .C(address_c_0), 
         .D(address_c_3), .Z(n20756)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(49[33:40])
    defparam i15233_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_4_lut_adj_855 (.A(n15362), .B(n33910), .C(n33946), 
         .D(address_c_3), .Z(n33)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(49[33:40])
    defparam i1_2_lut_3_lut_4_lut_adj_855.init = 16'hfffe;
    LUT4 i24334_2_lut_rep_606 (.A(address_c_2), .B(address_c_4), .Z(n33910)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24334_2_lut_rep_606.init = 16'heeee;
    LUT4 i2_2_lut_rep_557_3_lut (.A(address_c_2), .B(address_c_4), .C(n15362), 
         .Z(n33861)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_2_lut_rep_557_3_lut.init = 16'hfefe;
    LUT4 i2_3_lut_rep_609 (.A(aes_core_ctrl_new_1__N_858[1]), .B(enc_ctrl_new_2__N_1045), 
         .C(encdec_reg), .Z(n33913)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i2_3_lut_rep_609.init = 16'h8080;
    LUT4 i1_2_lut_4_lut_adj_856 (.A(aes_core_ctrl_new_1__N_858[1]), .B(enc_ctrl_new_2__N_1045), 
         .C(encdec_reg), .D(n33915), .Z(round_ctr_we_adj_9437)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_2_lut_4_lut_adj_856.init = 16'hff80;
    LUT4 i25797_then_3_lut (.A(result_reg[76]), .B(address_c_1), .C(result_reg[12]), 
         .Z(n34005)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i25797_then_3_lut.init = 16'he2e2;
    LUT4 i25860_then_3_lut (.A(result_reg[35]), .B(address_c_0), .C(result_reg[3]), 
         .Z(n34047)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i25860_then_3_lut.init = 16'he2e2;
    LUT4 i25860_else_3_lut (.A(result_reg[99]), .B(address_c_0), .C(result_reg[67]), 
         .Z(n34046)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i25860_else_3_lut.init = 16'he2e2;
    LUT4 i25797_else_3_lut (.A(result_reg[108]), .B(address_c_1), .C(result_reg[44]), 
         .Z(n34004)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i25797_else_3_lut.init = 16'he2e2;
    LUT4 i1_2_lut_rep_635 (.A(cs_c), .B(we_c), .Z(n33939)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(46[33:35])
    defparam i1_2_lut_rep_635.init = 16'h8888;
    LUT4 i1_2_lut_rep_553_3_lut (.A(cs_c), .B(we_c), .C(address_c_3), 
         .Z(n33857)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(46[33:35])
    defparam i1_2_lut_rep_553_3_lut.init = 16'h0808;
    LUT4 equal_135_i3_2_lut_rep_636 (.A(address_c_0), .B(address_c_1), .Z(n33940)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(209[13:38])
    defparam equal_135_i3_2_lut_rep_636.init = 16'hdddd;
    LUT4 i27861_2_lut_2_lut_3_lut_4_lut (.A(address_c_0), .B(address_c_1), 
         .C(n33850), .D(address_c_2), .Z(clk_c_enable_355)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(209[13:38])
    defparam i27861_2_lut_2_lut_3_lut_4_lut.init = 16'h0020;
    LUT4 i27863_2_lut_3_lut_3_lut_4_lut (.A(address_c_0), .B(address_c_1), 
         .C(address_c_2), .D(n33850), .Z(clk_c_enable_227)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(209[13:38])
    defparam i27863_2_lut_3_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i14325_2_lut_rep_637 (.A(address_c_0), .B(address_c_1), .Z(n33941)) /* synthesis lut_function=(A (B)) */ ;
    defparam i14325_2_lut_rep_637.init = 16'h8888;
    LUT4 i27888_2_lut_2_lut_3_lut_4_lut (.A(address_c_0), .B(address_c_1), 
         .C(n33850), .D(address_c_2), .Z(clk_c_enable_291)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i27888_2_lut_2_lut_3_lut_4_lut.init = 16'h0080;
    LUT4 i2_2_lut_3_lut_4_lut (.A(address_c_0), .B(address_c_1), .C(n33850), 
         .D(address_c_2), .Z(clk_c_enable_163)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i2_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_638 (.A(dec_ctrl_new_2__N_2032), .B(aes_core_ctrl_new_1__N_858[1]), 
         .Z(n33942)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_2_lut_rep_638.init = 16'h8888;
    LUT4 i1_2_lut_rep_554_3_lut (.A(dec_ctrl_new_2__N_2032), .B(aes_core_ctrl_new_1__N_858[1]), 
         .C(encdec_reg), .Z(n33858)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_2_lut_rep_554_3_lut.init = 16'h0808;
    LUT4 i1_2_lut_3_lut_4_lut_adj_857 (.A(dec_ctrl_new_2__N_2032), .B(aes_core_ctrl_new_1__N_858[1]), 
         .C(n149), .D(encdec_reg), .Z(round_ctr_we)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_2_lut_3_lut_4_lut_adj_857.init = 16'hf0f8;
    LUT4 i25800_then_3_lut (.A(result_reg[77]), .B(address_c_1), .C(result_reg[13]), 
         .Z(n34008)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i25800_then_3_lut.init = 16'he2e2;
    LUT4 i25800_else_3_lut (.A(result_reg[109]), .B(address_c_1), .C(result_reg[45]), 
         .Z(n34007)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i25800_else_3_lut.init = 16'he2e2;
    LUT4 i7590_1_lut (.A(write_data_c_1), .Z(n13203)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(50[33:43])
    defparam i7590_1_lut.init = 16'h5555;
    LUT4 i1_4_lut_adj_858 (.A(n33861), .B(n33939), .C(n33949), .D(address_c_3), 
         .Z(n10461)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(46[33:35])
    defparam i1_4_lut_adj_858.init = 16'h0400;
    LUT4 i7589_1_lut (.A(write_data_c_0), .Z(n13202)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(50[33:43])
    defparam i7589_1_lut.init = 16'h5555;
    VLO i1 (.Z(GND_net));
    TSALL TSALL_INST (.TSALL(GND_net));
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    LUT4 i25803_then_3_lut (.A(result_reg[78]), .B(address_c_1), .C(result_reg[14]), 
         .Z(n34011)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i25803_then_3_lut.init = 16'he2e2;
    LUT4 i25803_else_3_lut (.A(result_reg[110]), .B(address_c_1), .C(result_reg[46]), 
         .Z(n34010)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i25803_else_3_lut.init = 16'he2e2;
    LUT4 i25809_then_3_lut (.A(result_reg[80]), .B(address_c_1), .C(result_reg[16]), 
         .Z(n34014)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i25809_then_3_lut.init = 16'he2e2;
    LUT4 i25809_else_3_lut (.A(result_reg[112]), .B(address_c_1), .C(result_reg[48]), 
         .Z(n34013)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i25809_else_3_lut.init = 16'he2e2;
    LUT4 i25812_then_3_lut (.A(result_reg[81]), .B(address_c_1), .C(result_reg[17]), 
         .Z(n34017)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i25812_then_3_lut.init = 16'he2e2;
    LUT4 i25812_else_3_lut (.A(result_reg[113]), .B(address_c_1), .C(result_reg[49]), 
         .Z(n34016)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i25812_else_3_lut.init = 16'he2e2;
    LUT4 i1_3_lut_4_lut_4_lut (.A(\key_mem_ctrl.num_rounds [2]), .B(n15484), 
         .C(\key_reg[3] [2]), .D(n33860), .Z(prev_key1_new_127__N_4787[2])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_859 (.A(\key_mem_ctrl.num_rounds [2]), .B(n17229), 
         .C(\key_reg[2] [31]), .D(n33860), .Z(prev_key1_new_127__N_4787[63])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_859.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_860 (.A(\key_mem_ctrl.num_rounds [2]), .B(n15424), 
         .C(\key_reg[3] [1]), .D(n33860), .Z(prev_key1_new_127__N_4787[1])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_860.init = 16'hccdc;
    LUT4 i26973_3_lut_3_lut (.A(\key_mem_ctrl.num_rounds [2]), .B(n152), 
         .C(n14930), .Z(n14934)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i26973_3_lut_3_lut.init = 16'he4e4;
    LUT4 i1_3_lut_4_lut_4_lut_adj_861 (.A(\key_mem_ctrl.num_rounds [2]), .B(n15544), 
         .C(\key_reg[3] [3]), .D(n33860), .Z(prev_key1_new_127__N_4787[3])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_861.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_862 (.A(\key_mem_ctrl.num_rounds [2]), .B(n15604), 
         .C(\key_reg[3] [4]), .D(n33860), .Z(prev_key1_new_127__N_4787[4])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_862.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_863 (.A(\key_mem_ctrl.num_rounds [2]), .B(n15664), 
         .C(\key_reg[3] [5]), .D(n33860), .Z(prev_key1_new_127__N_4787[5])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_863.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_864 (.A(\key_mem_ctrl.num_rounds [2]), .B(n15724), 
         .C(\key_reg[3] [6]), .D(n33860), .Z(prev_key1_new_127__N_4787[6])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_864.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_865 (.A(\key_mem_ctrl.num_rounds [2]), .B(n15784), 
         .C(\key_reg[3] [7]), .D(n33860), .Z(prev_key1_new_127__N_4787[7])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_865.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_866 (.A(\key_mem_ctrl.num_rounds [2]), .B(n15844), 
         .C(\key_reg[3] [8]), .D(n33860), .Z(prev_key1_new_127__N_4787[8])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_866.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_867 (.A(\key_mem_ctrl.num_rounds [2]), .B(n15904), 
         .C(\key_reg[3] [9]), .D(n33860), .Z(prev_key1_new_127__N_4787[9])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_867.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_868 (.A(\key_mem_ctrl.num_rounds [2]), .B(n15964), 
         .C(\key_reg[3] [10]), .D(n33860), .Z(prev_key1_new_127__N_4787[10])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_868.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_869 (.A(\key_mem_ctrl.num_rounds [2]), .B(n16024), 
         .C(\key_reg[3] [11]), .D(n33860), .Z(prev_key1_new_127__N_4787[11])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_869.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_870 (.A(\key_mem_ctrl.num_rounds [2]), .B(n16084), 
         .C(\key_reg[3] [12]), .D(n33860), .Z(prev_key1_new_127__N_4787[12])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_870.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_871 (.A(\key_mem_ctrl.num_rounds [2]), .B(n16144), 
         .C(\key_reg[3] [13]), .D(n33860), .Z(prev_key1_new_127__N_4787[13])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_871.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_872 (.A(\key_mem_ctrl.num_rounds [2]), .B(n16204), 
         .C(\key_reg[3] [14]), .D(n33860), .Z(prev_key1_new_127__N_4787[14])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_872.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_873 (.A(\key_mem_ctrl.num_rounds [2]), .B(n16264), 
         .C(\key_reg[3] [15]), .D(n33860), .Z(prev_key1_new_127__N_4787[15])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_873.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_874 (.A(\key_mem_ctrl.num_rounds [2]), .B(n16324), 
         .C(\key_reg[3] [16]), .D(n33860), .Z(prev_key1_new_127__N_4787[16])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_874.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_875 (.A(\key_mem_ctrl.num_rounds [2]), .B(n16384), 
         .C(\key_reg[3] [17]), .D(n33860), .Z(prev_key1_new_127__N_4787[17])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_875.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_876 (.A(\key_mem_ctrl.num_rounds [2]), .B(n16444), 
         .C(\key_reg[3] [18]), .D(n33860), .Z(prev_key1_new_127__N_4787[18])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_876.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_877 (.A(\key_mem_ctrl.num_rounds [2]), .B(n16504), 
         .C(\key_reg[3] [19]), .D(n33860), .Z(prev_key1_new_127__N_4787[19])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_877.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_878 (.A(\key_mem_ctrl.num_rounds [2]), .B(n16564), 
         .C(\key_reg[3] [20]), .D(n33860), .Z(prev_key1_new_127__N_4787[20])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_878.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_879 (.A(\key_mem_ctrl.num_rounds [2]), .B(n16624), 
         .C(\key_reg[3] [21]), .D(n33860), .Z(prev_key1_new_127__N_4787[21])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_879.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_880 (.A(\key_mem_ctrl.num_rounds [2]), .B(n16684), 
         .C(\key_reg[3] [22]), .D(n33860), .Z(prev_key1_new_127__N_4787[22])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_880.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_881 (.A(\key_mem_ctrl.num_rounds [2]), .B(n16744), 
         .C(\key_reg[3] [23]), .D(n33860), .Z(prev_key1_new_127__N_4787[23])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_881.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_882 (.A(\key_mem_ctrl.num_rounds [2]), .B(n16804), 
         .C(\key_reg[3] [24]), .D(n33860), .Z(prev_key1_new_127__N_4787[24])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_882.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_883 (.A(\key_mem_ctrl.num_rounds [2]), .B(n16864), 
         .C(\key_reg[3] [25]), .D(n33860), .Z(prev_key1_new_127__N_4787[25])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_883.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_884 (.A(\key_mem_ctrl.num_rounds [2]), .B(n16924), 
         .C(\key_reg[3] [26]), .D(n33860), .Z(prev_key1_new_127__N_4787[26])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_884.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_885 (.A(\key_mem_ctrl.num_rounds [2]), .B(n16984), 
         .C(\key_reg[3] [27]), .D(n33860), .Z(prev_key1_new_127__N_4787[27])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_885.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_886 (.A(\key_mem_ctrl.num_rounds [2]), .B(n17044), 
         .C(\key_reg[3] [28]), .D(n33860), .Z(prev_key1_new_127__N_4787[28])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_886.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_887 (.A(\key_mem_ctrl.num_rounds [2]), .B(n17104), 
         .C(\key_reg[3] [29]), .D(n33860), .Z(prev_key1_new_127__N_4787[29])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_887.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_888 (.A(\key_mem_ctrl.num_rounds [2]), .B(n17164), 
         .C(\key_reg[3] [30]), .D(n33860), .Z(prev_key1_new_127__N_4787[30])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_888.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_889 (.A(\key_mem_ctrl.num_rounds [2]), .B(n17224), 
         .C(\key_reg[3] [31]), .D(n33860), .Z(prev_key1_new_127__N_4787[31])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_889.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_890 (.A(\key_mem_ctrl.num_rounds [2]), .B(n15316), 
         .C(\key_reg[2] [0]), .D(n33860), .Z(prev_key1_new_127__N_4787[32])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_890.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_891 (.A(\key_mem_ctrl.num_rounds [2]), .B(n15429), 
         .C(\key_reg[2] [1]), .D(n33860), .Z(prev_key1_new_127__N_4787[33])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_891.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_892 (.A(\key_mem_ctrl.num_rounds [2]), .B(n15489), 
         .C(\key_reg[2] [2]), .D(n33860), .Z(prev_key1_new_127__N_4787[34])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_892.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_893 (.A(\key_mem_ctrl.num_rounds [2]), .B(n15549), 
         .C(\key_reg[2] [3]), .D(n33860), .Z(prev_key1_new_127__N_4787[35])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_893.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_894 (.A(\key_mem_ctrl.num_rounds [2]), .B(n15609), 
         .C(\key_reg[2] [4]), .D(n33860), .Z(prev_key1_new_127__N_4787[36])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_894.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_895 (.A(\key_mem_ctrl.num_rounds [2]), .B(n15669), 
         .C(\key_reg[2] [5]), .D(n33860), .Z(prev_key1_new_127__N_4787[37])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_895.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_896 (.A(\key_mem_ctrl.num_rounds [2]), .B(n15729), 
         .C(\key_reg[2] [6]), .D(n33860), .Z(prev_key1_new_127__N_4787[38])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_896.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_897 (.A(\key_mem_ctrl.num_rounds [2]), .B(n15789), 
         .C(\key_reg[2] [7]), .D(n33860), .Z(prev_key1_new_127__N_4787[39])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_897.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_898 (.A(\key_mem_ctrl.num_rounds [2]), .B(n15849), 
         .C(\key_reg[2] [8]), .D(n33860), .Z(prev_key1_new_127__N_4787[40])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_898.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_899 (.A(\key_mem_ctrl.num_rounds [2]), .B(n15909), 
         .C(\key_reg[2] [9]), .D(n33860), .Z(prev_key1_new_127__N_4787[41])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_899.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_900 (.A(\key_mem_ctrl.num_rounds [2]), .B(n15969), 
         .C(\key_reg[2] [10]), .D(n33860), .Z(prev_key1_new_127__N_4787[42])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_900.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_901 (.A(\key_mem_ctrl.num_rounds [2]), .B(n16029), 
         .C(\key_reg[2] [11]), .D(n33860), .Z(prev_key1_new_127__N_4787[43])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_901.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_902 (.A(\key_mem_ctrl.num_rounds [2]), .B(n16089), 
         .C(\key_reg[2] [12]), .D(n33860), .Z(prev_key1_new_127__N_4787[44])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_902.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_903 (.A(\key_mem_ctrl.num_rounds [2]), .B(n16149), 
         .C(\key_reg[2] [13]), .D(n33860), .Z(prev_key1_new_127__N_4787[45])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_903.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_904 (.A(\key_mem_ctrl.num_rounds [2]), .B(n16209), 
         .C(\key_reg[2] [14]), .D(n33860), .Z(prev_key1_new_127__N_4787[46])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_904.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_905 (.A(\key_mem_ctrl.num_rounds [2]), .B(n16269), 
         .C(\key_reg[2] [15]), .D(n33860), .Z(prev_key1_new_127__N_4787[47])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_905.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_906 (.A(\key_mem_ctrl.num_rounds [2]), .B(n16329), 
         .C(\key_reg[2] [16]), .D(n33860), .Z(prev_key1_new_127__N_4787[48])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_906.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_907 (.A(\key_mem_ctrl.num_rounds [2]), .B(n16389), 
         .C(\key_reg[2] [17]), .D(n33860), .Z(prev_key1_new_127__N_4787[49])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_907.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_908 (.A(\key_mem_ctrl.num_rounds [2]), .B(n16449), 
         .C(\key_reg[2] [18]), .D(n33860), .Z(prev_key1_new_127__N_4787[50])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_908.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_909 (.A(\key_mem_ctrl.num_rounds [2]), .B(n16509), 
         .C(\key_reg[2] [19]), .D(n33860), .Z(prev_key1_new_127__N_4787[51])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_909.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_910 (.A(\key_mem_ctrl.num_rounds [2]), .B(n16569), 
         .C(\key_reg[2] [20]), .D(n33860), .Z(prev_key1_new_127__N_4787[52])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_910.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_911 (.A(\key_mem_ctrl.num_rounds [2]), .B(n16629), 
         .C(\key_reg[2] [21]), .D(n33860), .Z(prev_key1_new_127__N_4787[53])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_911.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_912 (.A(\key_mem_ctrl.num_rounds [2]), .B(n16689), 
         .C(\key_reg[2] [22]), .D(n33860), .Z(prev_key1_new_127__N_4787[54])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_912.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_913 (.A(\key_mem_ctrl.num_rounds [2]), .B(n16749), 
         .C(\key_reg[2] [23]), .D(n33860), .Z(prev_key1_new_127__N_4787[55])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_913.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_914 (.A(\key_mem_ctrl.num_rounds [2]), .B(n16809), 
         .C(\key_reg[2] [24]), .D(n33860), .Z(prev_key1_new_127__N_4787[56])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_914.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_915 (.A(\key_mem_ctrl.num_rounds [2]), .B(n16869), 
         .C(\key_reg[2] [25]), .D(n33860), .Z(prev_key1_new_127__N_4787[57])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_915.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_916 (.A(\key_mem_ctrl.num_rounds [2]), .B(n16929), 
         .C(\key_reg[2] [26]), .D(n33860), .Z(prev_key1_new_127__N_4787[58])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_916.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_917 (.A(\key_mem_ctrl.num_rounds [2]), .B(n16989), 
         .C(\key_reg[2] [27]), .D(n33860), .Z(prev_key1_new_127__N_4787[59])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_917.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_918 (.A(\key_mem_ctrl.num_rounds [2]), .B(n17049), 
         .C(\key_reg[2] [28]), .D(n33860), .Z(prev_key1_new_127__N_4787[60])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_918.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_919 (.A(\key_mem_ctrl.num_rounds [2]), .B(n17109), 
         .C(\key_reg[2] [29]), .D(n33860), .Z(prev_key1_new_127__N_4787[61])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_919.init = 16'hccdc;
    LUT4 i1_3_lut_4_lut_4_lut_adj_920 (.A(\key_mem_ctrl.num_rounds [2]), .B(n17169), 
         .C(\key_reg[2] [30]), .D(n33860), .Z(prev_key1_new_127__N_4787[62])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam i1_3_lut_4_lut_4_lut_adj_920.init = 16'hccdc;
    LUT4 address_7__I_0_111_i9_2_lut_rep_642 (.A(address_c_0), .B(address_c_1), 
         .Z(n33946)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(238[19:41])
    defparam address_7__I_0_111_i9_2_lut_rep_642.init = 16'hbbbb;
    LUT4 equal_42_i9_2_lut_rep_645 (.A(address_c_0), .B(address_c_1), .Z(n33949)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(251[17:27])
    defparam equal_42_i9_2_lut_rep_645.init = 16'heeee;
    LUT4 i1_2_lut_rep_646 (.A(we_c), .B(cs_c), .Z(n33950)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(46[33:35])
    defparam i1_2_lut_rep_646.init = 16'hbbbb;
    LUT4 i3417_2_lut_3_lut (.A(we_c), .B(cs_c), .C(n1504), .Z(n8904)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(46[33:35])
    defparam i3417_2_lut_3_lut.init = 16'h4040;
    LUT4 i25815_then_3_lut (.A(result_reg[82]), .B(address_c_1), .C(result_reg[18]), 
         .Z(n34020)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i25815_then_3_lut.init = 16'he2e2;
    LUT4 i25815_else_3_lut (.A(result_reg[114]), .B(address_c_1), .C(result_reg[50]), 
         .Z(n34019)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i25815_else_3_lut.init = 16'he2e2;
    LUT4 i25818_then_3_lut (.A(result_reg[83]), .B(address_c_1), .C(result_reg[19]), 
         .Z(n34023)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i25818_then_3_lut.init = 16'he2e2;
    LUT4 i25818_else_3_lut (.A(result_reg[115]), .B(address_c_1), .C(result_reg[51]), 
         .Z(n34022)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i25818_else_3_lut.init = 16'he2e2;
    LUT4 i25824_then_3_lut (.A(result_reg[85]), .B(address_c_1), .C(result_reg[21]), 
         .Z(n34026)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i25824_then_3_lut.init = 16'he2e2;
    LUT4 i25824_else_3_lut (.A(result_reg[117]), .B(address_c_1), .C(result_reg[53]), 
         .Z(n34025)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i25824_else_3_lut.init = 16'he2e2;
    LUT4 i25827_then_3_lut (.A(result_reg[86]), .B(address_c_1), .C(result_reg[22]), 
         .Z(n34029)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i25827_then_3_lut.init = 16'he2e2;
    LUT4 i25827_else_3_lut (.A(result_reg[118]), .B(address_c_1), .C(result_reg[54]), 
         .Z(n34028)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i25827_else_3_lut.init = 16'he2e2;
    LUT4 i1_3_lut (.A(address_c_5), .B(address_c_6), .C(address_c_7), 
         .Z(n28824)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;
    defparam i1_3_lut.init = 16'h0202;
    LUT4 i25833_then_3_lut (.A(result_reg[88]), .B(address_c_1), .C(result_reg[24]), 
         .Z(n34032)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i25833_then_3_lut.init = 16'he2e2;
    LUT4 i25833_else_3_lut (.A(result_reg[120]), .B(address_c_1), .C(result_reg[56]), 
         .Z(n34031)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i25833_else_3_lut.init = 16'he2e2;
    FD1P3AX keylen_reg_106_rep_650 (.D(write_data_c_1), .SP(config_we), 
            .CK(clk_c), .Q(n35835));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(192[9] 210[12])
    defparam keylen_reg_106_rep_650.GSR = "ENABLED";
    LUT4 i25845_then_3_lut (.A(result_reg[92]), .B(address_c_1), .C(result_reg[28]), 
         .Z(n34035)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i25845_then_3_lut.init = 16'he2e2;
    LUT4 i25845_else_3_lut (.A(result_reg[124]), .B(address_c_1), .C(result_reg[60]), 
         .Z(n34034)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i25845_else_3_lut.init = 16'he2e2;
    LUT4 i25848_then_3_lut (.A(result_reg[93]), .B(address_c_1), .C(result_reg[29]), 
         .Z(n34038)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i25848_then_3_lut.init = 16'he2e2;
    PFUMX i29020 (.BLUT(n33956), .ALUT(n33957), .C0(address_c_1), .Z(read_data_c_11));
    LUT4 i25848_else_3_lut (.A(result_reg[125]), .B(address_c_1), .C(result_reg[61]), 
         .Z(n34037)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i25848_else_3_lut.init = 16'he2e2;
    LUT4 i25851_then_3_lut (.A(result_reg[94]), .B(address_c_1), .C(result_reg[30]), 
         .Z(n34041)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i25851_then_3_lut.init = 16'he2e2;
    LUT4 i25851_else_3_lut (.A(result_reg[126]), .B(address_c_1), .C(result_reg[62]), 
         .Z(n34040)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i25851_else_3_lut.init = 16'he2e2;
    LUT4 i25857_then_3_lut (.A(result_reg[34]), .B(address_c_0), .C(result_reg[2]), 
         .Z(n34044)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i25857_then_3_lut.init = 16'he2e2;
    LUT4 i25857_else_3_lut (.A(result_reg[98]), .B(address_c_0), .C(result_reg[66]), 
         .Z(n34043)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i25857_else_3_lut.init = 16'he2e2;
    PFUMX i29080 (.BLUT(n34046), .ALUT(n34047), .C0(address_c_1), .Z(n34048));
    PFUMX i29018 (.BLUT(n33953), .ALUT(n33954), .C0(address_c_1), .Z(read_data_c_20));
    aes_core core (.encdec_reg(encdec_reg), .core_result({core_result}), 
            .\dec_round_nr[0] (dec_round_nr[0]), .aes_core_ctrl_reg({aes_core_ctrl_reg}), 
            .n33948(n33948), .core_ready(core_ready), .clk_c(clk_c), .ready_we(ready_we), 
            .core_valid(core_valid), .result_valid_we(result_valid_we), 
            .result_valid_new(result_valid_new), .n33947(n33947), .\key_mem_ctrl_new_2__N_4928[0] (key_mem_ctrl_new_2__N_4928[0]), 
            .\aes_core_ctrl_new_1__N_858[1] (aes_core_ctrl_new_1__N_858[1]), 
            .n1(n1), .n33860(n33860), .\key_reg[0] ({\key_reg[0] }), .n35835(n35835), 
            .GND_net(GND_net), .\new_sboxw[23] (new_sboxw[23]), .\new_sboxw[22] (new_sboxw[22]), 
            .\key_mem_ctrl.num_rounds[2] (\key_mem_ctrl.num_rounds [2]), .\key_reg[3] ({\key_reg[3] }), 
            .\key_reg[2] ({\key_reg[2] }), .\key_reg[1] ({\key_reg[1] }), 
            .\new_sboxw[21] (new_sboxw[21]), .\key_reg[5] ({\key_reg[5] }), 
            .\new_sboxw[20] (new_sboxw[20]), .\new_sboxw[19] (new_sboxw[19]), 
            .n15316(n15316), .\key_reg[6] ({\key_reg[6] }), .n15429(n15429), 
            .n15489(n15489), .n15549(n15549), .n15609(n15609), .n15669(n15669), 
            .n15729(n15729), .n15789(n15789), .n15849(n15849), .n15909(n15909), 
            .n15969(n15969), .n16029(n16029), .\new_sboxw[18] (new_sboxw[18]), 
            .\new_sboxw[17] (new_sboxw[17]), .n16089(n16089), .n16149(n16149), 
            .n16209(n16209), .n16269(n16269), .n16329(n16329), .\new_sboxw[16] (new_sboxw[16]), 
            .n16389(n16389), .n16449(n16449), .n16509(n16509), .n16569(n16569), 
            .n16629(n16629), .n16689(n16689), .n16749(n16749), .n16809(n16809), 
            .n16869(n16869), .n16929(n16929), .n16989(n16989), .n17049(n17049), 
            .n17109(n17109), .n17169(n17169), .n17229(n17229), .\key_reg[4] ({\key_reg[4] }), 
            .init_state(init_state), .\muxed_sboxw[16] (muxed_sboxw[16]), 
            .\muxed_sboxw[17] (muxed_sboxw[17]), .\muxed_sboxw[18] (muxed_sboxw[18]), 
            .\muxed_sboxw[19] (muxed_sboxw[19]), .\muxed_sboxw[20] (muxed_sboxw[20]), 
            .\muxed_sboxw[21] (muxed_sboxw[21]), .\muxed_sboxw[22] (muxed_sboxw[22]), 
            .\muxed_sboxw[23] (muxed_sboxw[23]), .reset_n_c(reset_n_c), 
            .\key_reg[7] ({\key_reg[7] }), .n17224(n17224), .n17164(n17164), 
            .n17104(n17104), .n17044(n17044), .n16984(n16984), .n16924(n16924), 
            .n16864(n16864), .n16804(n16804), .n16744(n16744), .n16684(n16684), 
            .n16624(n16624), .n16564(n16564), .n16504(n16504), .n16444(n16444), 
            .n16384(n16384), .n16324(n16324), .n16264(n16264), .n16204(n16204), 
            .n16144(n16144), .n16084(n16084), .n16024(n16024), .n15964(n15964), 
            .n15904(n15904), .n15844(n15844), .n15784(n15784), .n15724(n15724), 
            .n15664(n15664), .n15604(n15604), .n15544(n15544), .n15484(n15484), 
            .n15424(n15424), .\prev_key1_new_127__N_4787[1] (prev_key1_new_127__N_4787[1]), 
            .\prev_key1_new_127__N_4787[2] (prev_key1_new_127__N_4787[2]), 
            .\prev_key1_new_127__N_4787[3] (prev_key1_new_127__N_4787[3]), 
            .\prev_key1_new_127__N_4787[4] (prev_key1_new_127__N_4787[4]), 
            .\prev_key1_new_127__N_4787[5] (prev_key1_new_127__N_4787[5]), 
            .\prev_key1_new_127__N_4787[6] (prev_key1_new_127__N_4787[6]), 
            .\prev_key1_new_127__N_4787[7] (prev_key1_new_127__N_4787[7]), 
            .\prev_key1_new_127__N_4787[8] (prev_key1_new_127__N_4787[8]), 
            .\prev_key1_new_127__N_4787[9] (prev_key1_new_127__N_4787[9]), 
            .\prev_key1_new_127__N_4787[10] (prev_key1_new_127__N_4787[10]), 
            .\prev_key1_new_127__N_4787[11] (prev_key1_new_127__N_4787[11]), 
            .\prev_key1_new_127__N_4787[12] (prev_key1_new_127__N_4787[12]), 
            .\prev_key1_new_127__N_4787[13] (prev_key1_new_127__N_4787[13]), 
            .\prev_key1_new_127__N_4787[14] (prev_key1_new_127__N_4787[14]), 
            .\prev_key1_new_127__N_4787[15] (prev_key1_new_127__N_4787[15]), 
            .\prev_key1_new_127__N_4787[16] (prev_key1_new_127__N_4787[16]), 
            .\prev_key1_new_127__N_4787[17] (prev_key1_new_127__N_4787[17]), 
            .\prev_key1_new_127__N_4787[18] (prev_key1_new_127__N_4787[18]), 
            .\prev_key1_new_127__N_4787[19] (prev_key1_new_127__N_4787[19]), 
            .\prev_key1_new_127__N_4787[20] (prev_key1_new_127__N_4787[20]), 
            .\prev_key1_new_127__N_4787[21] (prev_key1_new_127__N_4787[21]), 
            .\prev_key1_new_127__N_4787[22] (prev_key1_new_127__N_4787[22]), 
            .\prev_key1_new_127__N_4787[23] (prev_key1_new_127__N_4787[23]), 
            .\prev_key1_new_127__N_4787[24] (prev_key1_new_127__N_4787[24]), 
            .\prev_key1_new_127__N_4787[25] (prev_key1_new_127__N_4787[25]), 
            .\prev_key1_new_127__N_4787[26] (prev_key1_new_127__N_4787[26]), 
            .\prev_key1_new_127__N_4787[27] (prev_key1_new_127__N_4787[27]), 
            .\prev_key1_new_127__N_4787[28] (prev_key1_new_127__N_4787[28]), 
            .\prev_key1_new_127__N_4787[29] (prev_key1_new_127__N_4787[29]), 
            .\prev_key1_new_127__N_4787[30] (prev_key1_new_127__N_4787[30]), 
            .\prev_key1_new_127__N_4787[31] (prev_key1_new_127__N_4787[31]), 
            .\prev_key1_new_127__N_4787[32] (prev_key1_new_127__N_4787[32]), 
            .\prev_key1_new_127__N_4787[33] (prev_key1_new_127__N_4787[33]), 
            .\prev_key1_new_127__N_4787[34] (prev_key1_new_127__N_4787[34]), 
            .\prev_key1_new_127__N_4787[35] (prev_key1_new_127__N_4787[35]), 
            .\prev_key1_new_127__N_4787[36] (prev_key1_new_127__N_4787[36]), 
            .\prev_key1_new_127__N_4787[37] (prev_key1_new_127__N_4787[37]), 
            .\prev_key1_new_127__N_4787[38] (prev_key1_new_127__N_4787[38]), 
            .\prev_key1_new_127__N_4787[39] (prev_key1_new_127__N_4787[39]), 
            .\prev_key1_new_127__N_4787[40] (prev_key1_new_127__N_4787[40]), 
            .\prev_key1_new_127__N_4787[41] (prev_key1_new_127__N_4787[41]), 
            .\prev_key1_new_127__N_4787[42] (prev_key1_new_127__N_4787[42]), 
            .\prev_key1_new_127__N_4787[43] (prev_key1_new_127__N_4787[43]), 
            .\prev_key1_new_127__N_4787[44] (prev_key1_new_127__N_4787[44]), 
            .\prev_key1_new_127__N_4787[45] (prev_key1_new_127__N_4787[45]), 
            .\prev_key1_new_127__N_4787[46] (prev_key1_new_127__N_4787[46]), 
            .\prev_key1_new_127__N_4787[47] (prev_key1_new_127__N_4787[47]), 
            .\prev_key1_new_127__N_4787[48] (prev_key1_new_127__N_4787[48]), 
            .\prev_key1_new_127__N_4787[49] (prev_key1_new_127__N_4787[49]), 
            .\prev_key1_new_127__N_4787[50] (prev_key1_new_127__N_4787[50]), 
            .\prev_key1_new_127__N_4787[51] (prev_key1_new_127__N_4787[51]), 
            .\prev_key1_new_127__N_4787[52] (prev_key1_new_127__N_4787[52]), 
            .\prev_key1_new_127__N_4787[53] (prev_key1_new_127__N_4787[53]), 
            .\prev_key1_new_127__N_4787[54] (prev_key1_new_127__N_4787[54]), 
            .\prev_key1_new_127__N_4787[55] (prev_key1_new_127__N_4787[55]), 
            .\prev_key1_new_127__N_4787[56] (prev_key1_new_127__N_4787[56]), 
            .\prev_key1_new_127__N_4787[57] (prev_key1_new_127__N_4787[57]), 
            .\prev_key1_new_127__N_4787[58] (prev_key1_new_127__N_4787[58]), 
            .\prev_key1_new_127__N_4787[59] (prev_key1_new_127__N_4787[59]), 
            .\prev_key1_new_127__N_4787[60] (prev_key1_new_127__N_4787[60]), 
            .\prev_key1_new_127__N_4787[61] (prev_key1_new_127__N_4787[61]), 
            .\prev_key1_new_127__N_4787[62] (prev_key1_new_127__N_4787[62]), 
            .\prev_key1_new_127__N_4787[63] (prev_key1_new_127__N_4787[63]), 
            .\block_reg[0] ({\block_reg[0] }), .\block_reg[1] ({\block_reg[1] }), 
            .enc_ctrl_new_2__N_1045(enc_ctrl_new_2__N_1045), .\block_reg[2] ({\block_reg[2] }), 
            .n33913(n33913), .round_ctr_we(round_ctr_we_adj_9437), .n33915(n33915), 
            .\block_reg[3] ({\block_reg[3] }), .tmp_sboxw({tmp_sboxw}), 
            .round_ctr_we_adj_128(round_ctr_we), .\round_ctr_new[0] (round_ctr_new[0]), 
            .n33858(n33858), .n149(n149), .new_sboxw({new_sboxw_adj_9440}), 
            .dec_ctrl_we(dec_ctrl_we), .n14934(n14934), .dec_ctrl_new_2__N_2032(dec_ctrl_new_2__N_2032), 
            .\round_ctr_new[3] (round_ctr_new[3]), .n33942(n33942), .n14930(n14930), 
            .n33909(n33909), .n14939(n14939), .n152(n152)) /* synthesis syn_module_defined=1 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(146[12] 161[17])
    
endmodule
//
// Verilog Description of module TSALL
// module not written out since it is a black-box. 
//

//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

//
// Verilog Description of module aes_core
//

module aes_core (encdec_reg, core_result, \dec_round_nr[0] , aes_core_ctrl_reg, 
            n33948, core_ready, clk_c, ready_we, core_valid, result_valid_we, 
            result_valid_new, n33947, \key_mem_ctrl_new_2__N_4928[0] , 
            \aes_core_ctrl_new_1__N_858[1] , n1, n33860, \key_reg[0] , 
            n35835, GND_net, \new_sboxw[23] , \new_sboxw[22] , \key_mem_ctrl.num_rounds[2] , 
            \key_reg[3] , \key_reg[2] , \key_reg[1] , \new_sboxw[21] , 
            \key_reg[5] , \new_sboxw[20] , \new_sboxw[19] , n15316, 
            \key_reg[6] , n15429, n15489, n15549, n15609, n15669, 
            n15729, n15789, n15849, n15909, n15969, n16029, \new_sboxw[18] , 
            \new_sboxw[17] , n16089, n16149, n16209, n16269, n16329, 
            \new_sboxw[16] , n16389, n16449, n16509, n16569, n16629, 
            n16689, n16749, n16809, n16869, n16929, n16989, n17049, 
            n17109, n17169, n17229, \key_reg[4] , init_state, \muxed_sboxw[16] , 
            \muxed_sboxw[17] , \muxed_sboxw[18] , \muxed_sboxw[19] , \muxed_sboxw[20] , 
            \muxed_sboxw[21] , \muxed_sboxw[22] , \muxed_sboxw[23] , reset_n_c, 
            \key_reg[7] , n17224, n17164, n17104, n17044, n16984, 
            n16924, n16864, n16804, n16744, n16684, n16624, n16564, 
            n16504, n16444, n16384, n16324, n16264, n16204, n16144, 
            n16084, n16024, n15964, n15904, n15844, n15784, n15724, 
            n15664, n15604, n15544, n15484, n15424, \prev_key1_new_127__N_4787[1] , 
            \prev_key1_new_127__N_4787[2] , \prev_key1_new_127__N_4787[3] , 
            \prev_key1_new_127__N_4787[4] , \prev_key1_new_127__N_4787[5] , 
            \prev_key1_new_127__N_4787[6] , \prev_key1_new_127__N_4787[7] , 
            \prev_key1_new_127__N_4787[8] , \prev_key1_new_127__N_4787[9] , 
            \prev_key1_new_127__N_4787[10] , \prev_key1_new_127__N_4787[11] , 
            \prev_key1_new_127__N_4787[12] , \prev_key1_new_127__N_4787[13] , 
            \prev_key1_new_127__N_4787[14] , \prev_key1_new_127__N_4787[15] , 
            \prev_key1_new_127__N_4787[16] , \prev_key1_new_127__N_4787[17] , 
            \prev_key1_new_127__N_4787[18] , \prev_key1_new_127__N_4787[19] , 
            \prev_key1_new_127__N_4787[20] , \prev_key1_new_127__N_4787[21] , 
            \prev_key1_new_127__N_4787[22] , \prev_key1_new_127__N_4787[23] , 
            \prev_key1_new_127__N_4787[24] , \prev_key1_new_127__N_4787[25] , 
            \prev_key1_new_127__N_4787[26] , \prev_key1_new_127__N_4787[27] , 
            \prev_key1_new_127__N_4787[28] , \prev_key1_new_127__N_4787[29] , 
            \prev_key1_new_127__N_4787[30] , \prev_key1_new_127__N_4787[31] , 
            \prev_key1_new_127__N_4787[32] , \prev_key1_new_127__N_4787[33] , 
            \prev_key1_new_127__N_4787[34] , \prev_key1_new_127__N_4787[35] , 
            \prev_key1_new_127__N_4787[36] , \prev_key1_new_127__N_4787[37] , 
            \prev_key1_new_127__N_4787[38] , \prev_key1_new_127__N_4787[39] , 
            \prev_key1_new_127__N_4787[40] , \prev_key1_new_127__N_4787[41] , 
            \prev_key1_new_127__N_4787[42] , \prev_key1_new_127__N_4787[43] , 
            \prev_key1_new_127__N_4787[44] , \prev_key1_new_127__N_4787[45] , 
            \prev_key1_new_127__N_4787[46] , \prev_key1_new_127__N_4787[47] , 
            \prev_key1_new_127__N_4787[48] , \prev_key1_new_127__N_4787[49] , 
            \prev_key1_new_127__N_4787[50] , \prev_key1_new_127__N_4787[51] , 
            \prev_key1_new_127__N_4787[52] , \prev_key1_new_127__N_4787[53] , 
            \prev_key1_new_127__N_4787[54] , \prev_key1_new_127__N_4787[55] , 
            \prev_key1_new_127__N_4787[56] , \prev_key1_new_127__N_4787[57] , 
            \prev_key1_new_127__N_4787[58] , \prev_key1_new_127__N_4787[59] , 
            \prev_key1_new_127__N_4787[60] , \prev_key1_new_127__N_4787[61] , 
            \prev_key1_new_127__N_4787[62] , \prev_key1_new_127__N_4787[63] , 
            \block_reg[0] , \block_reg[1] , enc_ctrl_new_2__N_1045, \block_reg[2] , 
            n33913, round_ctr_we, n33915, \block_reg[3] , tmp_sboxw, 
            round_ctr_we_adj_128, \round_ctr_new[0] , n33858, n149, 
            new_sboxw, dec_ctrl_we, n14934, dec_ctrl_new_2__N_2032, 
            \round_ctr_new[3] , n33942, n14930, n33909, n14939, n152) /* synthesis syn_module_defined=1 */ ;
    input encdec_reg;
    output [127:0]core_result;
    output \dec_round_nr[0] ;
    output [1:0]aes_core_ctrl_reg;
    output n33948;
    output core_ready;
    input clk_c;
    input ready_we;
    output core_valid;
    input result_valid_we;
    input result_valid_new;
    output n33947;
    input \key_mem_ctrl_new_2__N_4928[0] ;
    input \aes_core_ctrl_new_1__N_858[1] ;
    output n1;
    output n33860;
    input [31:0]\key_reg[0] ;
    input n35835;
    input GND_net;
    input \new_sboxw[23] ;
    input \new_sboxw[22] ;
    input \key_mem_ctrl.num_rounds[2] ;
    input [31:0]\key_reg[3] ;
    input [31:0]\key_reg[2] ;
    input [31:0]\key_reg[1] ;
    input \new_sboxw[21] ;
    input [31:0]\key_reg[5] ;
    input \new_sboxw[20] ;
    input \new_sboxw[19] ;
    output n15316;
    input [31:0]\key_reg[6] ;
    output n15429;
    output n15489;
    output n15549;
    output n15609;
    output n15669;
    output n15729;
    output n15789;
    output n15849;
    output n15909;
    output n15969;
    output n16029;
    input \new_sboxw[18] ;
    input \new_sboxw[17] ;
    output n16089;
    output n16149;
    output n16209;
    output n16269;
    output n16329;
    input \new_sboxw[16] ;
    output n16389;
    output n16449;
    output n16509;
    output n16569;
    output n16629;
    output n16689;
    output n16749;
    output n16809;
    output n16869;
    output n16929;
    output n16989;
    output n17049;
    output n17109;
    output n17169;
    output n17229;
    input [31:0]\key_reg[4] ;
    input init_state;
    output \muxed_sboxw[16] ;
    output \muxed_sboxw[17] ;
    output \muxed_sboxw[18] ;
    output \muxed_sboxw[19] ;
    output \muxed_sboxw[20] ;
    output \muxed_sboxw[21] ;
    output \muxed_sboxw[22] ;
    output \muxed_sboxw[23] ;
    input reset_n_c;
    input [31:0]\key_reg[7] ;
    output n17224;
    output n17164;
    output n17104;
    output n17044;
    output n16984;
    output n16924;
    output n16864;
    output n16804;
    output n16744;
    output n16684;
    output n16624;
    output n16564;
    output n16504;
    output n16444;
    output n16384;
    output n16324;
    output n16264;
    output n16204;
    output n16144;
    output n16084;
    output n16024;
    output n15964;
    output n15904;
    output n15844;
    output n15784;
    output n15724;
    output n15664;
    output n15604;
    output n15544;
    output n15484;
    output n15424;
    input \prev_key1_new_127__N_4787[1] ;
    input \prev_key1_new_127__N_4787[2] ;
    input \prev_key1_new_127__N_4787[3] ;
    input \prev_key1_new_127__N_4787[4] ;
    input \prev_key1_new_127__N_4787[5] ;
    input \prev_key1_new_127__N_4787[6] ;
    input \prev_key1_new_127__N_4787[7] ;
    input \prev_key1_new_127__N_4787[8] ;
    input \prev_key1_new_127__N_4787[9] ;
    input \prev_key1_new_127__N_4787[10] ;
    input \prev_key1_new_127__N_4787[11] ;
    input \prev_key1_new_127__N_4787[12] ;
    input \prev_key1_new_127__N_4787[13] ;
    input \prev_key1_new_127__N_4787[14] ;
    input \prev_key1_new_127__N_4787[15] ;
    input \prev_key1_new_127__N_4787[16] ;
    input \prev_key1_new_127__N_4787[17] ;
    input \prev_key1_new_127__N_4787[18] ;
    input \prev_key1_new_127__N_4787[19] ;
    input \prev_key1_new_127__N_4787[20] ;
    input \prev_key1_new_127__N_4787[21] ;
    input \prev_key1_new_127__N_4787[22] ;
    input \prev_key1_new_127__N_4787[23] ;
    input \prev_key1_new_127__N_4787[24] ;
    input \prev_key1_new_127__N_4787[25] ;
    input \prev_key1_new_127__N_4787[26] ;
    input \prev_key1_new_127__N_4787[27] ;
    input \prev_key1_new_127__N_4787[28] ;
    input \prev_key1_new_127__N_4787[29] ;
    input \prev_key1_new_127__N_4787[30] ;
    input \prev_key1_new_127__N_4787[31] ;
    input \prev_key1_new_127__N_4787[32] ;
    input \prev_key1_new_127__N_4787[33] ;
    input \prev_key1_new_127__N_4787[34] ;
    input \prev_key1_new_127__N_4787[35] ;
    input \prev_key1_new_127__N_4787[36] ;
    input \prev_key1_new_127__N_4787[37] ;
    input \prev_key1_new_127__N_4787[38] ;
    input \prev_key1_new_127__N_4787[39] ;
    input \prev_key1_new_127__N_4787[40] ;
    input \prev_key1_new_127__N_4787[41] ;
    input \prev_key1_new_127__N_4787[42] ;
    input \prev_key1_new_127__N_4787[43] ;
    input \prev_key1_new_127__N_4787[44] ;
    input \prev_key1_new_127__N_4787[45] ;
    input \prev_key1_new_127__N_4787[46] ;
    input \prev_key1_new_127__N_4787[47] ;
    input \prev_key1_new_127__N_4787[48] ;
    input \prev_key1_new_127__N_4787[49] ;
    input \prev_key1_new_127__N_4787[50] ;
    input \prev_key1_new_127__N_4787[51] ;
    input \prev_key1_new_127__N_4787[52] ;
    input \prev_key1_new_127__N_4787[53] ;
    input \prev_key1_new_127__N_4787[54] ;
    input \prev_key1_new_127__N_4787[55] ;
    input \prev_key1_new_127__N_4787[56] ;
    input \prev_key1_new_127__N_4787[57] ;
    input \prev_key1_new_127__N_4787[58] ;
    input \prev_key1_new_127__N_4787[59] ;
    input \prev_key1_new_127__N_4787[60] ;
    input \prev_key1_new_127__N_4787[61] ;
    input \prev_key1_new_127__N_4787[62] ;
    input \prev_key1_new_127__N_4787[63] ;
    input [31:0]\block_reg[0] ;
    input [31:0]\block_reg[1] ;
    output enc_ctrl_new_2__N_1045;
    input [31:0]\block_reg[2] ;
    input n33913;
    input round_ctr_we;
    output n33915;
    input [31:0]\block_reg[3] ;
    output [31:0]tmp_sboxw;
    input round_ctr_we_adj_128;
    input \round_ctr_new[0] ;
    input n33858;
    output n149;
    input [31:0]new_sboxw;
    input dec_ctrl_we;
    input n14934;
    output dec_ctrl_new_2__N_2032;
    input \round_ctr_new[3] ;
    input n33942;
    output n14930;
    output n33909;
    output n14939;
    output n152;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(41[33:36])
    wire [127:0]dec_new_block;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(100[18:31])
    wire [7:0]\round_logic.mixcolumns_block_7__N_1245 ;
    wire [127:0]enc_new_block;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(94[18:31])
    wire [7:0]\round_logic.mixcolumns_block_111__N_1285 ;
    wire [7:0]\round_logic.mixcolumns_block_39__N_1197 ;
    wire [7:0]\round_logic.mixcolumns_block_15__N_1453 ;
    wire [7:0]\round_logic.mixcolumns_block_71__N_1149 ;
    wire [7:0]\round_logic.mixcolumns_block_47__N_1397 ;
    wire [3:0]enc_round_nr;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(93[18:30])
    
    wire maxfan_replicated_net_23, key_ready, ready_new;
    wire [7:0]\round_logic.mixcolumns_block_79__N_1341 ;
    wire [7:0]\round_logic.mixcolumns_block_103__N_1101 ;
    
    wire n2634, n33952;
    wire [3:0]muxed_round_nr;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(104[18:32])
    
    wire n11;
    wire [127:0]\key_mem[14] ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(75[17:24])
    
    wire n33463, n11_adj_9293, n33462, n11_adj_9294, n33461, n11_adj_9295, 
        n33460, n11_adj_9296, n33459, n11_adj_9297, n33458, n11_adj_9298, 
        n33457, n11_adj_9299, n33456, n11_adj_9300, n33455, n11_adj_9301, 
        n33454, n11_adj_9302, n33453, n11_adj_9303, n33452, n11_adj_9304, 
        n33451, n11_adj_9305, n33450, n11_adj_9306, n33449, n11_adj_9307, 
        n33448, n11_adj_9308, n33447, n11_adj_9309, n33446, n11_adj_9310, 
        n33445, n11_adj_9311, n33444, n11_adj_9312, n33443, n11_adj_9313, 
        n33442, n11_adj_9314, n33441, n11_adj_9315, n33440, n11_adj_9316, 
        n33439, n11_adj_9317, n33438, n11_adj_9318, n33437, n11_adj_9319, 
        n33436, n11_adj_9320, n33435, n11_adj_9321, n33434, n11_adj_9322, 
        n33433, n11_adj_9323, n33432, n11_adj_9324, n33431, n11_adj_9325, 
        n33430, n11_adj_9326, n33429, n11_adj_9327, n33428, n11_adj_9328, 
        n33427, n11_adj_9329, n33426, n11_adj_9330, n33425, n11_adj_9331, 
        n33424, n11_adj_9332, n33423, n11_adj_9333, n33422, n11_adj_9334, 
        n33421, n11_adj_9335, n33420, n11_adj_9336, n33419, n11_adj_9337, 
        n33418, n11_adj_9338, n33417, n11_adj_9339, n33416, n11_adj_9340, 
        n33415, n11_adj_9341, n33414, n11_adj_9342, n33413, n11_adj_9343, 
        n33412, n11_adj_9344, n33411, n11_adj_9345, n33410, n11_adj_9346, 
        n33409, n11_adj_9347, n33408, n11_adj_9348, n33407, n11_adj_9349, 
        n33406, n11_adj_9350, n33405, n11_adj_9351, n33404, n11_adj_9352, 
        n33403, n11_adj_9353, n33402, n11_adj_9354, n33401, n11_adj_9355, 
        n33400, n11_adj_9356, n33399, n11_adj_9357, n33398, n11_adj_9358, 
        n33397, n11_adj_9359, n33396, n11_adj_9360, n33395, n11_adj_9361, 
        n33394, n11_adj_9362, n33393, n11_adj_9363, n33392, n11_adj_9364, 
        n33391, n11_adj_9365, n33390, n11_adj_9366, n33389, n11_adj_9367, 
        n33388, n11_adj_9368, n33387, n11_adj_9369, n33386, n11_adj_9370, 
        n33385, n11_adj_9371, n33384, n11_adj_9372, n33383, n11_adj_9373, 
        n33382, n11_adj_9374, n33381, n11_adj_9375, n33380, n11_adj_9376, 
        n33379, n11_adj_9377, n33378, n11_adj_9378, n33377, n11_adj_9379, 
        n33376, n11_adj_9380, n33375, n11_adj_9381, n33374, n11_adj_9382, 
        n33373, n11_adj_9383, n33372, n11_adj_9384, n33371, n11_adj_9385, 
        n33370, n11_adj_9386, n33369, n11_adj_9387, n33368, n11_adj_9388, 
        n33367, n11_adj_9389, n33366, n11_adj_9390, n33365, n11_adj_9391, 
        n33364, n11_adj_9392, n33363, n11_adj_9393, n33362, n11_adj_9394, 
        n33361, n11_adj_9395, n33360, n11_adj_9396, n33359, n11_adj_9397, 
        n33358, n11_adj_9398, n33357, n11_adj_9399, n33356, n11_adj_9400, 
        n33355, n11_adj_9401, n33354, n11_adj_9402, n33353, n11_adj_9403, 
        n33352, n11_adj_9404, n33351, n11_adj_9405, n33350, n11_adj_9406, 
        n33349, n11_adj_9407, n33348, n11_adj_9408, n33347, n11_adj_9409, 
        n33346, n11_adj_9410, n33345, n11_adj_9411, n33344, n11_adj_9412, 
        n33343, n11_adj_9413, n33342, n11_adj_9414, n33341, n11_adj_9415, 
        n33340, n11_adj_9416, n33339, n11_adj_9417, n33338, n11_adj_9418, 
        n33337, n11_adj_9419, n33336, dec_ready, enc_ready;
    wire [31:0]\round_key_gen.trw ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(191[39:42])
    
    wire n5;
    wire [127:0]round_key;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(89[18:27])
    wire [31:0]n2531;
    
    wire n8532, n9616, n9618, n9620, n9622, n9624, n9626, n9628, 
        n9630, n9632, n9634, n9636, n9638, n9640, n9642, n9644, 
        n9646, n9648, n9650, n9652, n9654, n9656, n9658, n9660, 
        n9662, n9664, n9666, n9668, n9670, n9672, n9674, n9676;
    wire [3:0]n6364;
    wire [3:0]n6347;
    
    wire n33846, n6428;
    wire [127:0]block_new_127__N_1645;
    
    wire n33848, n28773, n4;
    
    LUT4 dec_new_block_127__I_0_i38_3_lut (.A(dec_new_block[37]), .B(\round_logic.mixcolumns_block_7__N_1245 [6]), 
         .C(encdec_reg), .Z(core_result[37])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i38_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i39_3_lut (.A(dec_new_block[38]), .B(\round_logic.mixcolumns_block_7__N_1245 [7]), 
         .C(encdec_reg), .Z(core_result[38])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i39_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i40_3_lut (.A(dec_new_block[39]), .B(\round_logic.mixcolumns_block_7__N_1245 [0]), 
         .C(encdec_reg), .Z(core_result[39])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i40_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i41_3_lut (.A(dec_new_block[40]), .B(enc_new_block[40]), 
         .C(encdec_reg), .Z(core_result[40])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i41_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i42_3_lut (.A(dec_new_block[41]), .B(\round_logic.mixcolumns_block_111__N_1285 [2]), 
         .C(encdec_reg), .Z(core_result[41])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i42_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i43_3_lut (.A(dec_new_block[42]), .B(enc_new_block[42]), 
         .C(encdec_reg), .Z(core_result[42])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i43_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i44_3_lut (.A(dec_new_block[43]), .B(enc_new_block[43]), 
         .C(encdec_reg), .Z(core_result[43])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i44_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i45_3_lut (.A(dec_new_block[44]), .B(\round_logic.mixcolumns_block_111__N_1285 [5]), 
         .C(encdec_reg), .Z(core_result[44])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i45_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i46_3_lut (.A(dec_new_block[45]), .B(\round_logic.mixcolumns_block_111__N_1285 [6]), 
         .C(encdec_reg), .Z(core_result[45])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i46_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i47_3_lut (.A(dec_new_block[46]), .B(\round_logic.mixcolumns_block_111__N_1285 [7]), 
         .C(encdec_reg), .Z(core_result[46])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i47_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i48_3_lut (.A(dec_new_block[47]), .B(\round_logic.mixcolumns_block_111__N_1285 [0]), 
         .C(encdec_reg), .Z(core_result[47])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i48_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i49_3_lut (.A(dec_new_block[48]), .B(enc_new_block[48]), 
         .C(encdec_reg), .Z(core_result[48])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i49_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i50_3_lut (.A(dec_new_block[49]), .B(enc_new_block[49]), 
         .C(encdec_reg), .Z(core_result[49])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i50_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i51_3_lut (.A(dec_new_block[50]), .B(enc_new_block[50]), 
         .C(encdec_reg), .Z(core_result[50])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i51_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i52_3_lut (.A(dec_new_block[51]), .B(enc_new_block[51]), 
         .C(encdec_reg), .Z(core_result[51])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i52_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i53_3_lut (.A(dec_new_block[52]), .B(enc_new_block[52]), 
         .C(encdec_reg), .Z(core_result[52])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i53_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i54_3_lut (.A(dec_new_block[53]), .B(enc_new_block[53]), 
         .C(encdec_reg), .Z(core_result[53])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i54_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i55_3_lut (.A(dec_new_block[54]), .B(enc_new_block[54]), 
         .C(encdec_reg), .Z(core_result[54])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i55_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i56_3_lut (.A(dec_new_block[55]), .B(enc_new_block[55]), 
         .C(encdec_reg), .Z(core_result[55])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i56_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i57_3_lut (.A(dec_new_block[56]), .B(enc_new_block[56]), 
         .C(encdec_reg), .Z(core_result[56])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i57_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i58_3_lut (.A(dec_new_block[57]), .B(enc_new_block[57]), 
         .C(encdec_reg), .Z(core_result[57])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i58_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i59_3_lut (.A(dec_new_block[58]), .B(enc_new_block[58]), 
         .C(encdec_reg), .Z(core_result[58])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i59_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i60_3_lut (.A(dec_new_block[59]), .B(enc_new_block[59]), 
         .C(encdec_reg), .Z(core_result[59])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i60_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i61_3_lut (.A(dec_new_block[60]), .B(enc_new_block[60]), 
         .C(encdec_reg), .Z(core_result[60])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i61_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i62_3_lut (.A(dec_new_block[61]), .B(enc_new_block[61]), 
         .C(encdec_reg), .Z(core_result[61])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i62_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i63_3_lut (.A(dec_new_block[62]), .B(enc_new_block[62]), 
         .C(encdec_reg), .Z(core_result[62])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i63_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i64_3_lut (.A(dec_new_block[63]), .B(enc_new_block[63]), 
         .C(encdec_reg), .Z(core_result[63])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i64_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i65_3_lut (.A(dec_new_block[64]), .B(enc_new_block[64]), 
         .C(encdec_reg), .Z(core_result[64])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i65_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i66_3_lut (.A(dec_new_block[65]), .B(\round_logic.mixcolumns_block_39__N_1197 [2]), 
         .C(encdec_reg), .Z(core_result[65])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i66_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i67_3_lut (.A(dec_new_block[66]), .B(enc_new_block[66]), 
         .C(encdec_reg), .Z(core_result[66])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i67_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i68_3_lut (.A(dec_new_block[67]), .B(enc_new_block[67]), 
         .C(encdec_reg), .Z(core_result[67])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i68_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i69_3_lut (.A(dec_new_block[68]), .B(\round_logic.mixcolumns_block_39__N_1197 [5]), 
         .C(encdec_reg), .Z(core_result[68])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i69_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i70_3_lut (.A(dec_new_block[69]), .B(\round_logic.mixcolumns_block_39__N_1197 [6]), 
         .C(encdec_reg), .Z(core_result[69])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i70_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i71_3_lut (.A(dec_new_block[70]), .B(\round_logic.mixcolumns_block_39__N_1197 [7]), 
         .C(encdec_reg), .Z(core_result[70])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i71_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i72_3_lut (.A(dec_new_block[71]), .B(\round_logic.mixcolumns_block_39__N_1197 [0]), 
         .C(encdec_reg), .Z(core_result[71])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i72_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i73_3_lut (.A(dec_new_block[72]), .B(enc_new_block[72]), 
         .C(encdec_reg), .Z(core_result[72])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i73_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i74_3_lut (.A(dec_new_block[73]), .B(\round_logic.mixcolumns_block_15__N_1453 [2]), 
         .C(encdec_reg), .Z(core_result[73])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i74_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i75_3_lut (.A(dec_new_block[74]), .B(enc_new_block[74]), 
         .C(encdec_reg), .Z(core_result[74])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i75_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i76_3_lut (.A(dec_new_block[75]), .B(enc_new_block[75]), 
         .C(encdec_reg), .Z(core_result[75])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i76_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i77_3_lut (.A(dec_new_block[76]), .B(\round_logic.mixcolumns_block_15__N_1453 [5]), 
         .C(encdec_reg), .Z(core_result[76])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i77_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i78_3_lut (.A(dec_new_block[77]), .B(\round_logic.mixcolumns_block_15__N_1453 [6]), 
         .C(encdec_reg), .Z(core_result[77])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i78_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i79_3_lut (.A(dec_new_block[78]), .B(\round_logic.mixcolumns_block_15__N_1453 [7]), 
         .C(encdec_reg), .Z(core_result[78])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i79_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i80_3_lut (.A(dec_new_block[79]), .B(\round_logic.mixcolumns_block_15__N_1453 [0]), 
         .C(encdec_reg), .Z(core_result[79])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i80_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i81_3_lut (.A(dec_new_block[80]), .B(enc_new_block[80]), 
         .C(encdec_reg), .Z(core_result[80])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i81_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i82_3_lut (.A(dec_new_block[81]), .B(enc_new_block[81]), 
         .C(encdec_reg), .Z(core_result[81])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i82_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i83_3_lut (.A(dec_new_block[82]), .B(enc_new_block[82]), 
         .C(encdec_reg), .Z(core_result[82])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i83_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i84_3_lut (.A(dec_new_block[83]), .B(enc_new_block[83]), 
         .C(encdec_reg), .Z(core_result[83])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i84_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i85_3_lut (.A(dec_new_block[84]), .B(enc_new_block[84]), 
         .C(encdec_reg), .Z(core_result[84])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i85_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i86_3_lut (.A(dec_new_block[85]), .B(enc_new_block[85]), 
         .C(encdec_reg), .Z(core_result[85])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i86_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i87_3_lut (.A(dec_new_block[86]), .B(enc_new_block[86]), 
         .C(encdec_reg), .Z(core_result[86])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i87_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i88_3_lut (.A(dec_new_block[87]), .B(enc_new_block[87]), 
         .C(encdec_reg), .Z(core_result[87])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i88_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i89_3_lut (.A(dec_new_block[88]), .B(enc_new_block[88]), 
         .C(encdec_reg), .Z(core_result[88])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i89_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i90_3_lut (.A(dec_new_block[89]), .B(enc_new_block[89]), 
         .C(encdec_reg), .Z(core_result[89])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i90_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i91_3_lut (.A(dec_new_block[90]), .B(enc_new_block[90]), 
         .C(encdec_reg), .Z(core_result[90])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i91_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i92_3_lut (.A(dec_new_block[91]), .B(enc_new_block[91]), 
         .C(encdec_reg), .Z(core_result[91])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i92_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i93_3_lut (.A(dec_new_block[92]), .B(enc_new_block[92]), 
         .C(encdec_reg), .Z(core_result[92])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i93_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i94_3_lut (.A(dec_new_block[93]), .B(enc_new_block[93]), 
         .C(encdec_reg), .Z(core_result[93])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i94_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i95_3_lut (.A(dec_new_block[94]), .B(enc_new_block[94]), 
         .C(encdec_reg), .Z(core_result[94])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i95_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i96_3_lut (.A(dec_new_block[95]), .B(enc_new_block[95]), 
         .C(encdec_reg), .Z(core_result[95])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i96_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i97_3_lut (.A(dec_new_block[96]), .B(enc_new_block[96]), 
         .C(encdec_reg), .Z(core_result[96])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i97_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i98_3_lut (.A(dec_new_block[97]), .B(\round_logic.mixcolumns_block_71__N_1149 [2]), 
         .C(encdec_reg), .Z(core_result[97])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i98_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i99_3_lut (.A(dec_new_block[98]), .B(enc_new_block[98]), 
         .C(encdec_reg), .Z(core_result[98])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i99_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i100_3_lut (.A(dec_new_block[99]), .B(enc_new_block[99]), 
         .C(encdec_reg), .Z(core_result[99])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i100_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i101_3_lut (.A(dec_new_block[100]), .B(\round_logic.mixcolumns_block_71__N_1149 [5]), 
         .C(encdec_reg), .Z(core_result[100])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i101_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i102_3_lut (.A(dec_new_block[101]), .B(\round_logic.mixcolumns_block_71__N_1149 [6]), 
         .C(encdec_reg), .Z(core_result[101])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i102_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i103_3_lut (.A(dec_new_block[102]), .B(\round_logic.mixcolumns_block_71__N_1149 [7]), 
         .C(encdec_reg), .Z(core_result[102])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i103_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i104_3_lut (.A(dec_new_block[103]), .B(\round_logic.mixcolumns_block_71__N_1149 [0]), 
         .C(encdec_reg), .Z(core_result[103])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i104_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i105_3_lut (.A(dec_new_block[104]), .B(enc_new_block[104]), 
         .C(encdec_reg), .Z(core_result[104])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i105_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i106_3_lut (.A(dec_new_block[105]), .B(\round_logic.mixcolumns_block_47__N_1397 [2]), 
         .C(encdec_reg), .Z(core_result[105])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i106_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i107_3_lut (.A(dec_new_block[106]), .B(enc_new_block[106]), 
         .C(encdec_reg), .Z(core_result[106])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i107_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i108_3_lut (.A(dec_new_block[107]), .B(enc_new_block[107]), 
         .C(encdec_reg), .Z(core_result[107])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i108_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i109_3_lut (.A(dec_new_block[108]), .B(\round_logic.mixcolumns_block_47__N_1397 [5]), 
         .C(encdec_reg), .Z(core_result[108])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i109_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i110_3_lut (.A(dec_new_block[109]), .B(\round_logic.mixcolumns_block_47__N_1397 [6]), 
         .C(encdec_reg), .Z(core_result[109])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i110_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i111_3_lut (.A(dec_new_block[110]), .B(\round_logic.mixcolumns_block_47__N_1397 [7]), 
         .C(encdec_reg), .Z(core_result[110])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i111_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i112_3_lut (.A(dec_new_block[111]), .B(\round_logic.mixcolumns_block_47__N_1397 [0]), 
         .C(encdec_reg), .Z(core_result[111])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i112_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i113_3_lut (.A(dec_new_block[112]), .B(enc_new_block[112]), 
         .C(encdec_reg), .Z(core_result[112])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i113_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i114_3_lut (.A(dec_new_block[113]), .B(enc_new_block[113]), 
         .C(encdec_reg), .Z(core_result[113])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i114_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i115_3_lut (.A(dec_new_block[114]), .B(enc_new_block[114]), 
         .C(encdec_reg), .Z(core_result[114])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i115_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i116_3_lut (.A(dec_new_block[115]), .B(enc_new_block[115]), 
         .C(encdec_reg), .Z(core_result[115])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i116_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i117_3_lut (.A(dec_new_block[116]), .B(enc_new_block[116]), 
         .C(encdec_reg), .Z(core_result[116])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i117_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i118_3_lut (.A(dec_new_block[117]), .B(enc_new_block[117]), 
         .C(encdec_reg), .Z(core_result[117])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i118_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i119_3_lut (.A(dec_new_block[118]), .B(enc_new_block[118]), 
         .C(encdec_reg), .Z(core_result[118])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i119_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i120_3_lut (.A(dec_new_block[119]), .B(enc_new_block[119]), 
         .C(encdec_reg), .Z(core_result[119])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i120_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i121_3_lut (.A(dec_new_block[120]), .B(enc_new_block[120]), 
         .C(encdec_reg), .Z(core_result[120])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i121_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i122_3_lut (.A(dec_new_block[121]), .B(enc_new_block[121]), 
         .C(encdec_reg), .Z(core_result[121])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i122_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i123_3_lut (.A(dec_new_block[122]), .B(enc_new_block[122]), 
         .C(encdec_reg), .Z(core_result[122])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i123_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i124_3_lut (.A(dec_new_block[123]), .B(enc_new_block[123]), 
         .C(encdec_reg), .Z(core_result[123])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i124_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i125_3_lut (.A(dec_new_block[124]), .B(enc_new_block[124]), 
         .C(encdec_reg), .Z(core_result[124])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i125_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i126_3_lut (.A(dec_new_block[125]), .B(enc_new_block[125]), 
         .C(encdec_reg), .Z(core_result[125])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i126_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i127_3_lut (.A(dec_new_block[126]), .B(enc_new_block[126]), 
         .C(encdec_reg), .Z(core_result[126])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i127_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i128_3_lut (.A(dec_new_block[127]), .B(enc_new_block[127]), 
         .C(encdec_reg), .Z(core_result[127])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i128_3_lut.init = 16'hcaca;
    LUT4 dec_round_nr_3__I_0_i1_3_lut_rep_696 (.A(\dec_round_nr[0] ), .B(enc_round_nr[0]), 
         .C(encdec_reg), .Z(maxfan_replicated_net_23)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_round_nr_3__I_0_i1_3_lut_rep_696.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i27_3_lut (.A(dec_new_block[26]), .B(enc_new_block[26]), 
         .C(encdec_reg), .Z(core_result[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i27_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i26_3_lut (.A(dec_new_block[25]), .B(enc_new_block[25]), 
         .C(encdec_reg), .Z(core_result[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i26_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i25_3_lut (.A(dec_new_block[24]), .B(enc_new_block[24]), 
         .C(encdec_reg), .Z(core_result[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i25_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i24_3_lut (.A(dec_new_block[23]), .B(enc_new_block[23]), 
         .C(encdec_reg), .Z(core_result[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i24_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut (.A(aes_core_ctrl_reg[0]), .B(key_ready), .C(n33948), 
         .D(aes_core_ctrl_reg[1]), .Z(ready_new)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(195[9] 204[12])
    defparam i1_4_lut.init = 16'ha088;
    FD1P3AY ready_reg_32 (.D(ready_new), .SP(ready_we), .CK(clk_c), .Q(core_ready));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(195[9] 204[12])
    defparam ready_reg_32.GSR = "ENABLED";
    LUT4 dec_new_block_127__I_0_i28_3_lut (.A(dec_new_block[27]), .B(enc_new_block[27]), 
         .C(encdec_reg), .Z(core_result[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i28_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i23_3_lut (.A(dec_new_block[22]), .B(enc_new_block[22]), 
         .C(encdec_reg), .Z(core_result[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i23_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i29_3_lut (.A(dec_new_block[28]), .B(enc_new_block[28]), 
         .C(encdec_reg), .Z(core_result[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i29_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i30_3_lut (.A(dec_new_block[29]), .B(enc_new_block[29]), 
         .C(encdec_reg), .Z(core_result[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i30_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i31_3_lut (.A(dec_new_block[30]), .B(enc_new_block[30]), 
         .C(encdec_reg), .Z(core_result[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i31_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i32_3_lut (.A(dec_new_block[31]), .B(enc_new_block[31]), 
         .C(encdec_reg), .Z(core_result[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i32_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i33_3_lut (.A(dec_new_block[32]), .B(enc_new_block[32]), 
         .C(encdec_reg), .Z(core_result[32])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i33_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i34_3_lut (.A(dec_new_block[33]), .B(\round_logic.mixcolumns_block_7__N_1245 [2]), 
         .C(encdec_reg), .Z(core_result[33])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i34_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i35_3_lut (.A(dec_new_block[34]), .B(enc_new_block[34]), 
         .C(encdec_reg), .Z(core_result[34])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i35_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i36_3_lut (.A(dec_new_block[35]), .B(enc_new_block[35]), 
         .C(encdec_reg), .Z(core_result[35])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i36_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i37_3_lut (.A(dec_new_block[36]), .B(\round_logic.mixcolumns_block_7__N_1245 [5]), 
         .C(encdec_reg), .Z(core_result[36])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i37_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i22_3_lut (.A(dec_new_block[21]), .B(enc_new_block[21]), 
         .C(encdec_reg), .Z(core_result[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i22_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i21_3_lut (.A(dec_new_block[20]), .B(enc_new_block[20]), 
         .C(encdec_reg), .Z(core_result[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i21_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i20_3_lut (.A(dec_new_block[19]), .B(enc_new_block[19]), 
         .C(encdec_reg), .Z(core_result[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i20_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i19_3_lut (.A(dec_new_block[18]), .B(enc_new_block[18]), 
         .C(encdec_reg), .Z(core_result[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i19_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i18_3_lut (.A(dec_new_block[17]), .B(enc_new_block[17]), 
         .C(encdec_reg), .Z(core_result[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i18_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i1_3_lut (.A(dec_new_block[0]), .B(enc_new_block[0]), 
         .C(encdec_reg), .Z(core_result[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i1_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i17_3_lut (.A(dec_new_block[16]), .B(enc_new_block[16]), 
         .C(encdec_reg), .Z(core_result[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i17_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i16_3_lut (.A(dec_new_block[15]), .B(\round_logic.mixcolumns_block_79__N_1341 [0]), 
         .C(encdec_reg), .Z(core_result[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i16_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i15_3_lut (.A(dec_new_block[14]), .B(\round_logic.mixcolumns_block_79__N_1341 [7]), 
         .C(encdec_reg), .Z(core_result[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i15_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i14_3_lut (.A(dec_new_block[13]), .B(\round_logic.mixcolumns_block_79__N_1341 [6]), 
         .C(encdec_reg), .Z(core_result[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i14_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i13_3_lut (.A(dec_new_block[12]), .B(\round_logic.mixcolumns_block_79__N_1341 [5]), 
         .C(encdec_reg), .Z(core_result[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i13_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i12_3_lut (.A(dec_new_block[11]), .B(enc_new_block[11]), 
         .C(encdec_reg), .Z(core_result[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i12_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i11_3_lut (.A(dec_new_block[10]), .B(enc_new_block[10]), 
         .C(encdec_reg), .Z(core_result[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i11_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i10_3_lut (.A(dec_new_block[9]), .B(\round_logic.mixcolumns_block_79__N_1341 [2]), 
         .C(encdec_reg), .Z(core_result[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i10_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i9_3_lut (.A(dec_new_block[8]), .B(enc_new_block[8]), 
         .C(encdec_reg), .Z(core_result[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i9_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i8_3_lut (.A(dec_new_block[7]), .B(\round_logic.mixcolumns_block_103__N_1101 [0]), 
         .C(encdec_reg), .Z(core_result[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i8_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i7_3_lut (.A(dec_new_block[6]), .B(\round_logic.mixcolumns_block_103__N_1101 [7]), 
         .C(encdec_reg), .Z(core_result[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i7_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i6_3_lut (.A(dec_new_block[5]), .B(\round_logic.mixcolumns_block_103__N_1101 [6]), 
         .C(encdec_reg), .Z(core_result[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i6_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i5_3_lut (.A(dec_new_block[4]), .B(\round_logic.mixcolumns_block_103__N_1101 [5]), 
         .C(encdec_reg), .Z(core_result[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i5_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i4_3_lut (.A(dec_new_block[3]), .B(enc_new_block[3]), 
         .C(encdec_reg), .Z(core_result[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i4_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i3_3_lut (.A(dec_new_block[2]), .B(enc_new_block[2]), 
         .C(encdec_reg), .Z(core_result[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i3_3_lut.init = 16'hcaca;
    LUT4 dec_new_block_127__I_0_i2_3_lut (.A(dec_new_block[1]), .B(\round_logic.mixcolumns_block_103__N_1101 [2]), 
         .C(encdec_reg), .Z(core_result[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_new_block_127__I_0_i2_3_lut.init = 16'hcaca;
    FD1P3AX result_valid_reg_30 (.D(result_valid_new), .SP(result_valid_we), 
            .CK(clk_c), .Q(core_valid));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(195[9] 204[12])
    defparam result_valid_reg_30.GSR = "ENABLED";
    FD1P3IX aes_core_ctrl_reg_i0_i1 (.D(n2634), .SP(ready_we), .CD(ready_new), 
            .CK(clk_c), .Q(aes_core_ctrl_reg[1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=12, LSE_RCOL=17, LSE_LLINE=146, LSE_RLINE=161 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(195[9] 204[12])
    defparam aes_core_ctrl_reg_i0_i1.GSR = "ENABLED";
    FD1P3IX aes_core_ctrl_reg_i0_i0 (.D(n33947), .SP(ready_we), .CD(ready_new), 
            .CK(clk_c), .Q(aes_core_ctrl_reg[0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=12, LSE_RCOL=17, LSE_LLINE=146, LSE_RLINE=161 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(195[9] 204[12])
    defparam aes_core_ctrl_reg_i0_i0.GSR = "ENABLED";
    LUT4 \key_mem_14[[103__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11), .D(\key_mem[14] [103]), .Z(n33463)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[103__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[102__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9293), .D(\key_mem[14] [102]), .Z(n33462)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[102__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[101__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9294), .D(\key_mem[14] [101]), .Z(n33461)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[101__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[100__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9295), .D(\key_mem[14] [100]), .Z(n33460)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[100__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[99__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9296), .D(\key_mem[14] [99]), .Z(n33459)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[99__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[98__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9297), .D(\key_mem[14] [98]), .Z(n33458)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[98__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[97__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9298), .D(\key_mem[14] [97]), .Z(n33457)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[97__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[96__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9299), .D(\key_mem[14] [96]), .Z(n33456)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[96__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[95__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9300), .D(\key_mem[14] [95]), .Z(n33455)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[95__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[94__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9301), .D(\key_mem[14] [94]), .Z(n33454)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[94__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[93__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9302), .D(\key_mem[14] [93]), .Z(n33453)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[93__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[92__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9303), .D(\key_mem[14] [92]), .Z(n33452)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[92__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[91__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9304), .D(\key_mem[14] [91]), .Z(n33451)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[91__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[90__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9305), .D(\key_mem[14] [90]), .Z(n33450)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[90__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[89__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9306), .D(\key_mem[14] [89]), .Z(n33449)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[89__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[88__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9307), .D(\key_mem[14] [88]), .Z(n33448)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[88__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[114__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9308), .D(\key_mem[14] [114]), .Z(n33447)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[114__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[87__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9309), .D(\key_mem[14] [87]), .Z(n33446)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[87__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[113__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9310), .D(\key_mem[14] [113]), .Z(n33445)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[113__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[112__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9311), .D(\key_mem[14] [112]), .Z(n33444)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[112__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[111__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9312), .D(\key_mem[14] [111]), .Z(n33443)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[111__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[110__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9313), .D(\key_mem[14] [110]), .Z(n33442)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[110__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[86__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9314), .D(\key_mem[14] [86]), .Z(n33441)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[86__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[109__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9315), .D(\key_mem[14] [109]), .Z(n33440)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[109__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[108__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9316), .D(\key_mem[14] [108]), .Z(n33439)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[108__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[107__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9317), .D(\key_mem[14] [107]), .Z(n33438)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[107__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[106__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9318), .D(\key_mem[14] [106]), .Z(n33437)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[106__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[85__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9319), .D(\key_mem[14] [85]), .Z(n33436)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[85__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[105__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9320), .D(\key_mem[14] [105]), .Z(n33435)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[105__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[84__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9321), .D(\key_mem[14] [84]), .Z(n33434)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[84__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[83__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9322), .D(\key_mem[14] [83]), .Z(n33433)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[83__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[82__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9323), .D(\key_mem[14] [82]), .Z(n33432)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[82__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[81__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9324), .D(\key_mem[14] [81]), .Z(n33431)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[81__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[80__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9325), .D(\key_mem[14] [80]), .Z(n33430)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[80__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[79__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9326), .D(\key_mem[14] [79]), .Z(n33429)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[79__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[78__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9327), .D(\key_mem[14] [78]), .Z(n33428)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[78__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[77__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9328), .D(\key_mem[14] [77]), .Z(n33427)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[77__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[76__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9329), .D(\key_mem[14] [76]), .Z(n33426)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[76__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[75__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9330), .D(\key_mem[14] [75]), .Z(n33425)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[75__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[74__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9331), .D(\key_mem[14] [74]), .Z(n33424)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[74__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[73__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9332), .D(\key_mem[14] [73]), .Z(n33423)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[73__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[72__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9333), .D(\key_mem[14] [72]), .Z(n33422)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[72__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[71__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9334), .D(\key_mem[14] [71]), .Z(n33421)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[71__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[70__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9335), .D(\key_mem[14] [70]), .Z(n33420)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[70__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[69__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9336), .D(\key_mem[14] [69]), .Z(n33419)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[69__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[68__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9337), .D(\key_mem[14] [68]), .Z(n33418)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[68__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[67__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9338), .D(\key_mem[14] [67]), .Z(n33417)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[67__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[66__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9339), .D(\key_mem[14] [66]), .Z(n33416)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[66__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[65__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9340), .D(\key_mem[14] [65]), .Z(n33415)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[65__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[64__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9341), .D(\key_mem[14] [64]), .Z(n33414)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[64__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[42__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9342), .D(\key_mem[14] [42]), .Z(n33413)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[42__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[63__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9343), .D(\key_mem[14] [63]), .Z(n33412)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[63__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[41__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9344), .D(\key_mem[14] [41]), .Z(n33411)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[41__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[62__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9345), .D(\key_mem[14] [62]), .Z(n33410)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[62__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[40__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9346), .D(\key_mem[14] [40]), .Z(n33409)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[40__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[61__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9347), .D(\key_mem[14] [61]), .Z(n33408)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[61__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[60__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9348), .D(\key_mem[14] [60]), .Z(n33407)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[60__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[39__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9349), .D(\key_mem[14] [39]), .Z(n33406)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[39__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[38__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9350), .D(\key_mem[14] [38]), .Z(n33405)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[38__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[59__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9351), .D(\key_mem[14] [59]), .Z(n33404)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[59__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[58__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9352), .D(\key_mem[14] [58]), .Z(n33403)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[58__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[37__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9353), .D(\key_mem[14] [37]), .Z(n33402)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[37__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[57__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9354), .D(\key_mem[14] [57]), .Z(n33401)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[57__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[36__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9355), .D(\key_mem[14] [36]), .Z(n33400)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[36__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[56__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9356), .D(\key_mem[14] [56]), .Z(n33399)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[56__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[35__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9357), .D(\key_mem[14] [35]), .Z(n33398)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[35__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[55__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9358), .D(\key_mem[14] [55]), .Z(n33397)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[55__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[54__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9359), .D(\key_mem[14] [54]), .Z(n33396)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[54__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[34__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9360), .D(\key_mem[14] [34]), .Z(n33395)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[34__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[53__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9361), .D(\key_mem[14] [53]), .Z(n33394)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[53__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[33__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9362), .D(\key_mem[14] [33]), .Z(n33393)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[33__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[52__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9363), .D(\key_mem[14] [52]), .Z(n33392)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[52__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[32__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9364), .D(\key_mem[14] [32]), .Z(n33391)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[32__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[51__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9365), .D(\key_mem[14] [51]), .Z(n33390)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[51__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[31__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9366), .D(\key_mem[14] [31]), .Z(n33389)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[31__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[24__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9367), .D(\key_mem[14] [24]), .Z(n33388)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[24__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[30__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9368), .D(\key_mem[14] [30]), .Z(n33387)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[30__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[29__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9369), .D(\key_mem[14] [29]), .Z(n33386)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[29__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[23__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9370), .D(\key_mem[14] [23]), .Z(n33385)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[23__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[28__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9371), .D(\key_mem[14] [28]), .Z(n33384)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[28__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[22__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9372), .D(\key_mem[14] [22]), .Z(n33383)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[22__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[27__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9373), .D(\key_mem[14] [27]), .Z(n33382)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[27__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[21__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9374), .D(\key_mem[14] [21]), .Z(n33381)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[21__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[25__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9375), .D(\key_mem[14] [25]), .Z(n33380)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[25__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[127__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9376), .D(\key_mem[14] [127]), .Z(n33379)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[127__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[20__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9377), .D(\key_mem[14] [20]), .Z(n33378)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[20__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[126__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9378), .D(\key_mem[14] [126]), .Z(n33377)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[126__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[50__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9379), .D(\key_mem[14] [50]), .Z(n33376)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[50__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[19__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9380), .D(\key_mem[14] [19]), .Z(n33375)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[19__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[125__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9381), .D(\key_mem[14] [125]), .Z(n33374)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[125__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[18__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9382), .D(\key_mem[14] [18]), .Z(n33373)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[18__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[17__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9383), .D(\key_mem[14] [17]), .Z(n33372)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[17__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[49__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9384), .D(\key_mem[14] [49]), .Z(n33371)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[49__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[48__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9385), .D(\key_mem[14] [48]), .Z(n33370)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[48__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[47__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9386), .D(\key_mem[14] [47]), .Z(n33369)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[47__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[16__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9387), .D(\key_mem[14] [16]), .Z(n33368)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[16__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[124__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9388), .D(\key_mem[14] [124]), .Z(n33367)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[124__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[15__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9389), .D(\key_mem[14] [15]), .Z(n33366)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[15__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[14__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9390), .D(\key_mem[14] [14]), .Z(n33365)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[14__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[13__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9391), .D(\key_mem[14] [13]), .Z(n33364)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[13__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[12__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9392), .D(\key_mem[14] [12]), .Z(n33363)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[12__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[11__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9393), .D(\key_mem[14] [11]), .Z(n33362)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[11__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[123__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9394), .D(\key_mem[14] [123]), .Z(n33361)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[123__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[10__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9395), .D(\key_mem[14] [10]), .Z(n33360)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[10__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[9__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9396), .D(\key_mem[14] [9]), .Z(n33359)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[9__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[0__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9397), .D(\key_mem[14] [0]), .Z(n33358)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[0__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[8__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9398), .D(\key_mem[14] [8]), .Z(n33357)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[8__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[7__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9399), .D(\key_mem[14] [7]), .Z(n33356)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[7__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[122__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9400), .D(\key_mem[14] [122]), .Z(n33355)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[122__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[26__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9401), .D(\key_mem[14] [26]), .Z(n33354)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[26__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[6__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9402), .D(\key_mem[14] [6]), .Z(n33353)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[6__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[5__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9403), .D(\key_mem[14] [5]), .Z(n33352)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[5__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[4__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9404), .D(\key_mem[14] [4]), .Z(n33351)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[4__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[121__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9405), .D(\key_mem[14] [121]), .Z(n33350)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[121__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[3__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9406), .D(\key_mem[14] [3]), .Z(n33349)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[3__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[2__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9407), .D(\key_mem[14] [2]), .Z(n33348)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[2__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[1__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9408), .D(\key_mem[14] [1]), .Z(n33347)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[1__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[46__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9409), .D(\key_mem[14] [46]), .Z(n33346)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[46__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[45__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9410), .D(\key_mem[14] [45]), .Z(n33345)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[45__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[44__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9411), .D(\key_mem[14] [44]), .Z(n33344)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[44__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[43__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9412), .D(\key_mem[14] [43]), .Z(n33343)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[43__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[120__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9413), .D(\key_mem[14] [120]), .Z(n33342)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[120__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[119__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9414), .D(\key_mem[14] [119]), .Z(n33341)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[119__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[118__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9415), .D(\key_mem[14] [118]), .Z(n33340)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[118__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[117__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9416), .D(\key_mem[14] [117]), .Z(n33339)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[117__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[116__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9417), .D(\key_mem[14] [116]), .Z(n33338)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[116__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[115__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9418), .D(\key_mem[14] [115]), .Z(n33337)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[115__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 \key_mem_14[[104__bdd_4_lut_4_lut  (.A(n33952), .B(muxed_round_nr[1]), 
         .C(n11_adj_9419), .D(\key_mem[14] [104]), .Z(n33336)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam \key_mem_14[[104__bdd_4_lut_4_lut .init = 16'h7430;
    LUT4 i186_2_lut (.A(\key_mem_ctrl_new_2__N_4928[0] ), .B(\aes_core_ctrl_new_1__N_858[1] ), 
         .Z(n2634)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(287[18] 296[18])
    defparam i186_2_lut.init = 16'h4444;
    LUT4 i200_2_lut_rep_643 (.A(\key_mem_ctrl_new_2__N_4928[0] ), .B(\aes_core_ctrl_new_1__N_858[1] ), 
         .Z(n33947)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(274[7] 331[14])
    defparam i200_2_lut_rep_643.init = 16'heeee;
    LUT4 mux_194_Mux_0_i1_3_lut_4_lut (.A(\key_mem_ctrl_new_2__N_4928[0] ), 
         .B(\aes_core_ctrl_new_1__N_858[1] ), .C(aes_core_ctrl_reg[0]), 
         .D(key_ready), .Z(n1)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(274[7] 331[14])
    defparam mux_194_Mux_0_i1_3_lut_4_lut.init = 16'hfe0e;
    LUT4 i23_3_lut_rep_644 (.A(dec_ready), .B(enc_ready), .C(encdec_reg), 
         .Z(n33948)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(195[9] 204[12])
    defparam i23_3_lut_rep_644.init = 16'hcaca;
    LUT4 dec_round_nr_3__I_0_i1_3_lut_rep_648 (.A(\dec_round_nr[0] ), .B(enc_round_nr[0]), 
         .C(encdec_reg), .Z(n33952)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(247[9] 253[12])
    defparam dec_round_nr_3__I_0_i1_3_lut_rep_648.init = 16'hcaca;
    aes_key_mem keymem (.n33952(n33952), .\muxed_round_nr[1] (muxed_round_nr[1]), 
            .\round_key_gen.trw[2] (\round_key_gen.trw [2]), .n33860(n33860), 
            .\key_reg[0] ({\key_reg[0] }), .n11(n11_adj_9296), .\round_key_gen.trw[1] (\round_key_gen.trw [1]), 
            .n35835(n35835), .clk_c(clk_c), .GND_net(GND_net), .\round_key_gen.trw[0] (\round_key_gen.trw [0]), 
            .\new_sboxw[23] (\new_sboxw[23] ), .\new_sboxw[22] (\new_sboxw[22] ), 
            .\key_mem_ctrl.num_rounds[2] (\key_mem_ctrl.num_rounds[2] ), .\key_reg[3] ({\key_reg[3] }), 
            .\key_reg[2] ({\key_reg[2] }), .\key_reg[1] ({\key_reg[1] }), 
            .n11_adj_1(n11_adj_9297), .\new_sboxw[21] (\new_sboxw[21] ), 
            .\key_reg[5] ({\key_reg[5] }), .\new_sboxw[20] (\new_sboxw[20] ), 
            .\new_sboxw[19] (\new_sboxw[19] ), .n11_adj_2(n11_adj_9418), 
            .n11_adj_3(n11_adj_9308), .n15316(n15316), .\key_reg[6] ({\key_reg[6] }), 
            .\round_key_gen.trw[8] (\round_key_gen.trw [8]), .n15429(n15429), 
            .\round_key_gen.trw[9] (\round_key_gen.trw [9]), .n15489(n15489), 
            .\round_key_gen.trw[10] (\round_key_gen.trw [10]), .n15549(n15549), 
            .\round_key_gen.trw[3] (\round_key_gen.trw [3]), .\round_key_gen.trw[11] (\round_key_gen.trw [11]), 
            .n15609(n15609), .n11_adj_4(n11_adj_9309), .\round_key_gen.trw[4] (\round_key_gen.trw [4]), 
            .\round_key_gen.trw[12] (\round_key_gen.trw [12]), .n15669(n15669), 
            .\round_key_gen.trw[5] (\round_key_gen.trw [5]), .\round_key_gen.trw[13] (\round_key_gen.trw [13]), 
            .n15729(n15729), .\round_key_gen.trw[6] (\round_key_gen.trw [6]), 
            .\round_key_gen.trw[14] (\round_key_gen.trw [14]), .n15789(n15789), 
            .\round_key_gen.trw[7] (\round_key_gen.trw [7]), .\round_key_gen.trw[15] (\round_key_gen.trw [15]), 
            .n15849(n15849), .\round_key_gen.trw[16] (\round_key_gen.trw [16]), 
            .n11_adj_5(n11_adj_9298), .n15909(n15909), .n11_adj_6(n11_adj_9310), 
            .\round_key_gen.trw[17] (\round_key_gen.trw [17]), .n15969(n15969), 
            .\round_key_gen.trw[18] (\round_key_gen.trw [18]), .n16029(n16029), 
            .\new_sboxw[18] (\new_sboxw[18] ), .\round_key_gen.trw[19] (\round_key_gen.trw [19]), 
            .\new_sboxw[17] (\new_sboxw[17] ), .n11_adj_7(n11_adj_9311), 
            .n16089(n16089), .\round_key_gen.trw[20] (\round_key_gen.trw [20]), 
            .n16149(n16149), .\round_key_gen.trw[21] (\round_key_gen.trw [21]), 
            .n11_adj_8(n11_adj_9312), .n16209(n16209), .\round_key_gen.trw[22] (\round_key_gen.trw [22]), 
            .n16269(n16269), .\round_key_gen.trw[23] (\round_key_gen.trw [23]), 
            .n16329(n16329), .\new_sboxw[16] (\new_sboxw[16] ), .n11_adj_9(n11_adj_9313), 
            .n16389(n16389), .n11_adj_10(n11_adj_9314), .n16449(n16449), 
            .n11_adj_11(n11_adj_9315), .n16509(n16509), .n16569(n16569), 
            .n11_adj_12(n11_adj_9316), .n11_adj_13(n11_adj_9299), .n16629(n16629), 
            .n16689(n16689), .n11_adj_14(n11_adj_9317), .n16749(n16749), 
            .n16809(n16809), .n11_adj_15(n11_adj_9318), .n16869(n16869), 
            .n11_adj_16(n11_adj_9319), .n16929(n16929), .n11_adj_17(n11_adj_9320), 
            .n16989(n16989), .n17049(n17049), .n17109(n17109), .n17169(n17169), 
            .n11_adj_18(n11_adj_9321), .n17229(n17229), .n11_adj_19(n11_adj_9322), 
            .n11_adj_20(n11_adj_9323), .\key_reg[4] ({\key_reg[4] }), .n11_adj_21(n11_adj_9324), 
            .n11_adj_22(n11_adj_9325), .n11_adj_23(n11_adj_9300), .n11_adj_24(n11_adj_9326), 
            .n11_adj_25(n11_adj_9327), .n11_adj_26(n11_adj_9328), .n11_adj_27(n11_adj_9329), 
            .n11_adj_28(n11_adj_9330), .n11_adj_29(n11_adj_9331), .n11_adj_30(n11_adj_9332), 
            .n11_adj_31(n11_adj_9301), .n11_adj_32(n11_adj_9333), .n11_adj_33(n11_adj_9302), 
            .\key_mem[14] ({\key_mem[14] }), .n11_adj_34(n11_adj_9334), 
            .n5(n5), .init_state(init_state), .n11_adj_35(n11_adj_9335), 
            .n11_adj_36(n11_adj_9336), .n11_adj_37(n11_adj_9303), .n11_adj_38(n11_adj_9337), 
            .n11_adj_39(n11_adj_9338), .n11_adj_40(n11_adj_9304), .n11_adj_41(n11_adj_9339), 
            .\muxed_sboxw[16] (\muxed_sboxw[16] ), .\muxed_sboxw[17] (\muxed_sboxw[17] ), 
            .\muxed_sboxw[18] (\muxed_sboxw[18] ), .\muxed_sboxw[19] (\muxed_sboxw[19] ), 
            .\muxed_sboxw[20] (\muxed_sboxw[20] ), .n11_adj_42(n11_adj_9340), 
            .\muxed_sboxw[21] (\muxed_sboxw[21] ), .\muxed_sboxw[22] (\muxed_sboxw[22] ), 
            .\muxed_sboxw[23] (\muxed_sboxw[23] ), .key_ready(key_ready), 
            .n11_adj_43(n11_adj_9341), .n11_adj_44(n11_adj_9342), .n11_adj_45(n11_adj_9343), 
            .n11_adj_46(n11_adj_9344), .reset_n_c(reset_n_c), .n11_adj_47(n11_adj_9305), 
            .n11_adj_48(n11_adj_9306), .n11_adj_49(n11_adj_9307), .n11_adj_50(n11_adj_9345), 
            .n11_adj_51(n11_adj_9346), .n11_adj_52(n11_adj_9347), .n11_adj_53(n11_adj_9348), 
            .n11_adj_54(n11_adj_9349), .n11_adj_55(n11_adj_9350), .n11_adj_56(n11_adj_9351), 
            .n11_adj_57(n11_adj_9352), .n11_adj_58(n11_adj_9353), .n11_adj_59(n11_adj_9354), 
            .n11_adj_60(n11_adj_9355), .n11_adj_61(n11_adj_9356), .n11_adj_62(n11_adj_9357), 
            .n11_adj_63(n11_adj_9358), .n11_adj_64(n11_adj_9359), .n11_adj_65(n11_adj_9360), 
            .n11_adj_66(n11_adj_9361), .n11_adj_67(n11_adj_9362), .n11_adj_68(n11_adj_9363), 
            .n11_adj_69(n11_adj_9364), .n11_adj_70(n11_adj_9365), .n11_adj_71(n11_adj_9366), 
            .n11_adj_72(n11_adj_9367), .n11_adj_73(n11_adj_9368), .n11_adj_74(n11_adj_9369), 
            .n11_adj_75(n11_adj_9370), .n11_adj_76(n11_adj_9371), .n11_adj_77(n11_adj_9372), 
            .\muxed_round_nr[3] (muxed_round_nr[3]), .round_key({round_key}), 
            .n11_adj_78(n11_adj_9373), .n11_adj_79(n11_adj_9374), .n11_adj_80(n11_adj_9375), 
            .n11_adj_81(n11_adj_9376), .n11_adj_82(n11_adj_9377), .n11_adj_83(n11_adj_9378), 
            .n11_adj_84(n11_adj_9379), .n11_adj_85(n11_adj_9380), .n11_adj_86(n11_adj_9382), 
            .n11_adj_87(n11_adj_9381), .n11_adj_88(n11_adj_9383), .n11_adj_89(n11_adj_9384), 
            .\key_reg[7] ({\key_reg[7] }), .n11_adj_90(n11_adj_9385), .n11_adj_91(n11_adj_9386), 
            .n11_adj_92(n11_adj_9387), .n11_adj_93(n11_adj_9388), .n11_adj_94(n11_adj_9389), 
            .n11_adj_95(n11_adj_9390), .\muxed_round_nr[2] (muxed_round_nr[2]), 
            .n33343(n33343), .n33344(n33344), .n33345(n33345), .n33346(n33346), 
            .n33347(n33347), .n33348(n33348), .n33349(n33349), .n33351(n33351), 
            .n33352(n33352), .n33353(n33353), .n33354(n33354), .n33356(n33356), 
            .n33357(n33357), .n33358(n33358), .n33359(n33359), .n33360(n33360), 
            .n33362(n33362), .n33363(n33363), .n33364(n33364), .n33365(n33365), 
            .n11_adj_96(n11_adj_9391), .n33366(n33366), .n33368(n33368), 
            .n33369(n33369), .n33370(n33370), .n33371(n33371), .n11_adj_97(n11_adj_9392), 
            .n33372(n33372), .n33373(n33373), .n33375(n33375), .n33376(n33376), 
            .n33378(n33378), .n33381(n33381), .n33383(n33383), .n33385(n33385), 
            .n33388(n33388), .n33390(n33390), .n11_adj_98(n11_adj_9393), 
            .n11_adj_99(n11_adj_9395), .n11_adj_100(n11_adj_9394), .n33392(n33392), 
            .n11_adj_101(n11_adj_9396), .n17224(n17224), .n17164(n17164), 
            .n17104(n17104), .n11_adj_102(n11_adj_9397), .n17044(n17044), 
            .n16984(n16984), .n16924(n16924), .n16864(n16864), .n16804(n16804), 
            .n16744(n16744), .n16684(n16684), .n16624(n16624), .n11_adj_103(n11_adj_9398), 
            .n16564(n16564), .n16504(n16504), .n16444(n16444), .n16384(n16384), 
            .n16324(n16324), .n16264(n16264), .n16204(n16204), .n16144(n16144), 
            .n16084(n16084), .n11_adj_104(n11_adj_9399), .n16024(n16024), 
            .n15964(n15964), .n15904(n15904), .n15844(n15844), .n15784(n15784), 
            .n15724(n15724), .n15664(n15664), .n15604(n15604), .n15544(n15544), 
            .n15484(n15484), .n15424(n15424), .n11_adj_105(n11_adj_9400), 
            .n11_adj_106(n11_adj_9401), .n11_adj_107(n11_adj_9402), .n11_adj_108(n11_adj_9403), 
            .n11_adj_109(n11_adj_9404), .n11_adj_110(n11_adj_9405), .n11_adj_111(n11_adj_9406), 
            .n33394(n33394), .n11_adj_112(n11_adj_9407), .n33396(n33396), 
            .n33397(n33397), .n33399(n33399), .n33401(n33401), .n11_adj_113(n11_adj_9408), 
            .n33403(n33403), .n11_adj_114(n11_adj_9409), .maxfan_replicated_net_23(maxfan_replicated_net_23), 
            .n11_adj_115(n11_adj_9410), .n33404(n33404), .n33407(n33407), 
            .n33408(n33408), .n33410(n33410), .n11_adj_116(n11_adj_9411), 
            .n33412(n33412), .n33414(n33414), .n33415(n33415), .n33416(n33416), 
            .n11_adj_117(n11_adj_9412), .n33417(n33417), .n33418(n33418), 
            .n33419(n33419), .n33420(n33420), .n33421(n33421), .n33422(n33422), 
            .n33423(n33423), .n33424(n33424), .n33425(n33425), .n33426(n33426), 
            .n33427(n33427), .n33428(n33428), .n33429(n33429), .n33430(n33430), 
            .n11_adj_118(n11_adj_9413), .n11_adj_119(n11_adj_9414), .n11_adj_120(n11_adj_9415), 
            .n11_adj_121(n11_adj_9416), .n11_adj_122(n11_adj_9417), .\prev_key1_new_127__N_4787[1] (\prev_key1_new_127__N_4787[1] ), 
            .\prev_key1_new_127__N_4787[2] (\prev_key1_new_127__N_4787[2] ), 
            .\prev_key1_new_127__N_4787[3] (\prev_key1_new_127__N_4787[3] ), 
            .\prev_key1_new_127__N_4787[4] (\prev_key1_new_127__N_4787[4] ), 
            .\prev_key1_new_127__N_4787[5] (\prev_key1_new_127__N_4787[5] ), 
            .\prev_key1_new_127__N_4787[6] (\prev_key1_new_127__N_4787[6] ), 
            .\prev_key1_new_127__N_4787[7] (\prev_key1_new_127__N_4787[7] ), 
            .\prev_key1_new_127__N_4787[8] (\prev_key1_new_127__N_4787[8] ), 
            .\prev_key1_new_127__N_4787[9] (\prev_key1_new_127__N_4787[9] ), 
            .\prev_key1_new_127__N_4787[10] (\prev_key1_new_127__N_4787[10] ), 
            .\prev_key1_new_127__N_4787[11] (\prev_key1_new_127__N_4787[11] ), 
            .\prev_key1_new_127__N_4787[12] (\prev_key1_new_127__N_4787[12] ), 
            .\prev_key1_new_127__N_4787[13] (\prev_key1_new_127__N_4787[13] ), 
            .\prev_key1_new_127__N_4787[14] (\prev_key1_new_127__N_4787[14] ), 
            .\prev_key1_new_127__N_4787[15] (\prev_key1_new_127__N_4787[15] ), 
            .\prev_key1_new_127__N_4787[16] (\prev_key1_new_127__N_4787[16] ), 
            .\prev_key1_new_127__N_4787[17] (\prev_key1_new_127__N_4787[17] ), 
            .\prev_key1_new_127__N_4787[18] (\prev_key1_new_127__N_4787[18] ), 
            .\prev_key1_new_127__N_4787[19] (\prev_key1_new_127__N_4787[19] ), 
            .\prev_key1_new_127__N_4787[20] (\prev_key1_new_127__N_4787[20] ), 
            .\prev_key1_new_127__N_4787[21] (\prev_key1_new_127__N_4787[21] ), 
            .\prev_key1_new_127__N_4787[22] (\prev_key1_new_127__N_4787[22] ), 
            .\prev_key1_new_127__N_4787[23] (\prev_key1_new_127__N_4787[23] ), 
            .\prev_key1_new_127__N_4787[24] (\prev_key1_new_127__N_4787[24] ), 
            .\prev_key1_new_127__N_4787[25] (\prev_key1_new_127__N_4787[25] ), 
            .\prev_key1_new_127__N_4787[26] (\prev_key1_new_127__N_4787[26] ), 
            .\prev_key1_new_127__N_4787[27] (\prev_key1_new_127__N_4787[27] ), 
            .\prev_key1_new_127__N_4787[28] (\prev_key1_new_127__N_4787[28] ), 
            .\prev_key1_new_127__N_4787[29] (\prev_key1_new_127__N_4787[29] ), 
            .\prev_key1_new_127__N_4787[30] (\prev_key1_new_127__N_4787[30] ), 
            .\prev_key1_new_127__N_4787[31] (\prev_key1_new_127__N_4787[31] ), 
            .\prev_key1_new_127__N_4787[32] (\prev_key1_new_127__N_4787[32] ), 
            .\prev_key1_new_127__N_4787[33] (\prev_key1_new_127__N_4787[33] ), 
            .\prev_key1_new_127__N_4787[34] (\prev_key1_new_127__N_4787[34] ), 
            .\prev_key1_new_127__N_4787[35] (\prev_key1_new_127__N_4787[35] ), 
            .\prev_key1_new_127__N_4787[36] (\prev_key1_new_127__N_4787[36] ), 
            .\prev_key1_new_127__N_4787[37] (\prev_key1_new_127__N_4787[37] ), 
            .\prev_key1_new_127__N_4787[38] (\prev_key1_new_127__N_4787[38] ), 
            .\prev_key1_new_127__N_4787[39] (\prev_key1_new_127__N_4787[39] ), 
            .\prev_key1_new_127__N_4787[40] (\prev_key1_new_127__N_4787[40] ), 
            .\prev_key1_new_127__N_4787[41] (\prev_key1_new_127__N_4787[41] ), 
            .\prev_key1_new_127__N_4787[42] (\prev_key1_new_127__N_4787[42] ), 
            .\prev_key1_new_127__N_4787[43] (\prev_key1_new_127__N_4787[43] ), 
            .\prev_key1_new_127__N_4787[44] (\prev_key1_new_127__N_4787[44] ), 
            .\prev_key1_new_127__N_4787[45] (\prev_key1_new_127__N_4787[45] ), 
            .\prev_key1_new_127__N_4787[46] (\prev_key1_new_127__N_4787[46] ), 
            .\prev_key1_new_127__N_4787[47] (\prev_key1_new_127__N_4787[47] ), 
            .\prev_key1_new_127__N_4787[48] (\prev_key1_new_127__N_4787[48] ), 
            .\prev_key1_new_127__N_4787[49] (\prev_key1_new_127__N_4787[49] ), 
            .\prev_key1_new_127__N_4787[50] (\prev_key1_new_127__N_4787[50] ), 
            .\prev_key1_new_127__N_4787[51] (\prev_key1_new_127__N_4787[51] ), 
            .\prev_key1_new_127__N_4787[52] (\prev_key1_new_127__N_4787[52] ), 
            .\prev_key1_new_127__N_4787[53] (\prev_key1_new_127__N_4787[53] ), 
            .\prev_key1_new_127__N_4787[54] (\prev_key1_new_127__N_4787[54] ), 
            .\prev_key1_new_127__N_4787[55] (\prev_key1_new_127__N_4787[55] ), 
            .\prev_key1_new_127__N_4787[56] (\prev_key1_new_127__N_4787[56] ), 
            .\prev_key1_new_127__N_4787[57] (\prev_key1_new_127__N_4787[57] ), 
            .\prev_key1_new_127__N_4787[58] (\prev_key1_new_127__N_4787[58] ), 
            .\prev_key1_new_127__N_4787[59] (\prev_key1_new_127__N_4787[59] ), 
            .\prev_key1_new_127__N_4787[60] (\prev_key1_new_127__N_4787[60] ), 
            .\prev_key1_new_127__N_4787[61] (\prev_key1_new_127__N_4787[61] ), 
            .\prev_key1_new_127__N_4787[62] (\prev_key1_new_127__N_4787[62] ), 
            .\prev_key1_new_127__N_4787[63] (\prev_key1_new_127__N_4787[63] ), 
            .n33431(n33431), .n33432(n33432), .n11_adj_123(n11), .n33433(n33433), 
            .n33434(n33434), .n33436(n33436), .n33441(n33441), .n33446(n33446), 
            .n33448(n33448), .n33449(n33449), .n33450(n33450), .n33451(n33451), 
            .n33452(n33452), .n33453(n33453), .n33454(n33454), .n33455(n33455), 
            .n33456(n33456), .n33457(n33457), .n33458(n33458), .n33459(n33459), 
            .n33460(n33460), .n33461(n33461), .n11_adj_124(n11_adj_9293), 
            .n33462(n33462), .n33463(n33463), .n33336(n33336), .n33435(n33435), 
            .n33437(n33437), .n33438(n33438), .n33439(n33439), .n33440(n33440), 
            .n33442(n33442), .n33443(n33443), .n33444(n33444), .n33445(n33445), 
            .n33447(n33447), .n33337(n33337), .n33338(n33338), .n33339(n33339), 
            .n33340(n33340), .n33341(n33341), .n33342(n33342), .n33350(n33350), 
            .n33355(n33355), .n33361(n33361), .n33367(n33367), .n33374(n33374), 
            .n33377(n33377), .n33379(n33379), .n33380(n33380), .n33382(n33382), 
            .n33384(n33384), .n33386(n33386), .n11_adj_125(n11_adj_9294), 
            .n33387(n33387), .n33389(n33389), .n33391(n33391), .n33393(n33393), 
            .n33395(n33395), .n33398(n33398), .n33400(n33400), .n33402(n33402), 
            .n33405(n33405), .n33406(n33406), .n33409(n33409), .n33411(n33411), 
            .n33413(n33413), .n11_adj_126(n11_adj_9295), .n2531({n2531}), 
            .n8532(n8532), .n9616(n9616), .n9618(n9618), .n9620(n9620), 
            .n9622(n9622), .n9624(n9624), .n9626(n9626), .n9628(n9628), 
            .n9630(n9630), .n9632(n9632), .n9634(n9634), .n9636(n9636), 
            .n9638(n9638), .n9640(n9640), .n9642(n9642), .n9644(n9644), 
            .n9646(n9646), .n9648(n9648), .n9650(n9650), .n9652(n9652), 
            .n9654(n9654), .n9656(n9656), .n9658(n9658), .n9660(n9660), 
            .n9662(n9662), .n11_adj_127(n11_adj_9419), .n9664(n9664), 
            .n9666(n9666), .n9668(n9668), .n9670(n9670), .n9672(n9672), 
            .n9674(n9674), .n9676(n9676), .\key_mem_ctrl_new_2__N_4928[0] (\key_mem_ctrl_new_2__N_4928[0] ), 
            .block_w3_we_N_1490(n6364[3]), .block_w2_we_N_1489(n6364[2])) /* synthesis syn_module_defined=1 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(151[15] 165[22])
    aes_encipher_block enc_block (.n6347({enc_ctrl_new_2__N_1045, n6347[2:0]}), 
            .clk_c(clk_c), .\new_sboxw[19] (\new_sboxw[19] ), .n33846(n33846), 
            .\new_sboxw[20] (\new_sboxw[20] ), .enc_ready(enc_ready), .n6428(n6428), 
            .\new_sboxw[21] (\new_sboxw[21] ), .\round_key_gen.trw[1] (\round_key_gen.trw [1]), 
            .round_key({round_key}), .\block_reg[0][5] (\block_reg[0] [5]), 
            .\round_key_gen.trw[13] (\round_key_gen.trw [13]), .\block_reg[0][4] (\block_reg[0] [4]), 
            .\round_key_gen.trw[12] (\round_key_gen.trw [12]), .\block_reg[0][0] (\block_reg[0] [0]), 
            .\enc_new_block[56] (enc_new_block[56]), .\enc_new_block[24] (enc_new_block[24]), 
            .n6364({n6364[3], Open_0, Open_1, Open_2}), .n9662(n9662), 
            .\enc_new_block[120] (enc_new_block[120]), .\enc_new_block[88] (enc_new_block[88]), 
            .n2531({n2531}), .\enc_new_block[40] (enc_new_block[40]), .\round_key_gen.trw[8] (\round_key_gen.trw [8]), 
            .\block_reg[1][31] (\block_reg[1] [31]), .\round_key_gen.trw[3] (\round_key_gen.trw [3]), 
            .\enc_new_block[55] (enc_new_block[55]), .\enc_new_block[23] (enc_new_block[23]), 
            .n9660(n9660), .\enc_new_block[119] (enc_new_block[119]), .\enc_new_block[87] (enc_new_block[87]), 
            .\round_logic.mixcolumns_block_71__N_1149[0] (\round_logic.mixcolumns_block_71__N_1149 [0]), 
            .\round_key_gen.trw[7] (\round_key_gen.trw [7]), .\round_key_gen.trw[4] (\round_key_gen.trw [4]), 
            .\enc_new_block[54] (enc_new_block[54]), .\enc_new_block[22] (enc_new_block[22]), 
            .n9658(n9658), .\block_reg[1][30] (\block_reg[1] [30]), .\enc_new_block[118] (enc_new_block[118]), 
            .\enc_new_block[86] (enc_new_block[86]), .\round_key_gen.trw[6] (\round_key_gen.trw [6]), 
            .\enc_new_block[53] (enc_new_block[53]), .\enc_new_block[21] (enc_new_block[21]), 
            .n9656(n9656), .\enc_new_block[117] (enc_new_block[117]), .\enc_new_block[85] (enc_new_block[85]), 
            .\round_key_gen.trw[9] (\round_key_gen.trw [9]), .\round_key_gen.trw[10] (\round_key_gen.trw [10]), 
            .\enc_new_block[52] (enc_new_block[52]), .\enc_new_block[20] (enc_new_block[20]), 
            .n9654(n9654), .\block_reg[1][29] (\block_reg[1] [29]), .\enc_new_block[116] (enc_new_block[116]), 
            .\enc_new_block[84] (enc_new_block[84]), .\enc_new_block[51] (enc_new_block[51]), 
            .\enc_new_block[19] (enc_new_block[19]), .n9652(n9652), .\round_key_gen.trw[5] (\round_key_gen.trw [5]), 
            .\enc_new_block[115] (enc_new_block[115]), .\enc_new_block[83] (enc_new_block[83]), 
            .\round_key_gen.trw[11] (\round_key_gen.trw [11]), .\enc_new_block[50] (enc_new_block[50]), 
            .\enc_new_block[18] (enc_new_block[18]), .n9650(n9650), .\enc_new_block[58] (enc_new_block[58]), 
            .\round_key_gen.trw[14] (\round_key_gen.trw [14]), .\round_key_gen.trw[17] (\round_key_gen.trw [17]), 
            .\block_reg[1][26] (\block_reg[1] [26]), .\enc_new_block[114] (enc_new_block[114]), 
            .\enc_new_block[82] (enc_new_block[82]), .\round_key_gen.trw[19] (\round_key_gen.trw [19]), 
            .\enc_new_block[49] (enc_new_block[49]), .\enc_new_block[17] (enc_new_block[17]), 
            .n9648(n9648), .\enc_new_block[67] (enc_new_block[67]), .\enc_new_block[113] (enc_new_block[113]), 
            .\enc_new_block[81] (enc_new_block[81]), .\round_key_gen.trw[20] (\round_key_gen.trw [20]), 
            .\enc_new_block[48] (enc_new_block[48]), .\enc_new_block[16] (enc_new_block[16]), 
            .n9646(n9646), .\enc_new_block[112] (enc_new_block[112]), .\enc_new_block[80] (enc_new_block[80]), 
            .\round_logic.mixcolumns_block_111__N_1285[0] (\round_logic.mixcolumns_block_111__N_1285 [0]), 
            .\round_logic.mixcolumns_block_79__N_1341[0] (\round_logic.mixcolumns_block_79__N_1341 [0]), 
            .n9644(n9644), .\round_logic.mixcolumns_block_47__N_1397[0] (\round_logic.mixcolumns_block_47__N_1397 [0]), 
            .\round_logic.mixcolumns_block_15__N_1453[0] (\round_logic.mixcolumns_block_15__N_1453 [0]), 
            .\round_logic.mixcolumns_block_111__N_1285[7] (\round_logic.mixcolumns_block_111__N_1285 [7]), 
            .\round_logic.mixcolumns_block_79__N_1341[7] (\round_logic.mixcolumns_block_79__N_1341 [7]), 
            .n9642(n9642), .\round_logic.mixcolumns_block_47__N_1397[7] (\round_logic.mixcolumns_block_47__N_1397 [7]), 
            .\round_logic.mixcolumns_block_15__N_1453[7] (\round_logic.mixcolumns_block_15__N_1453 [7]), 
            .\new_sboxw[17] (\new_sboxw[17] ), .\round_logic.mixcolumns_block_111__N_1285[6] (\round_logic.mixcolumns_block_111__N_1285 [6]), 
            .\round_logic.mixcolumns_block_79__N_1341[6] (\round_logic.mixcolumns_block_79__N_1341 [6]), 
            .n9640(n9640), .\new_sboxw[18] (\new_sboxw[18] ), .\round_key_gen.trw[15] (\round_key_gen.trw [15]), 
            .\new_sboxw[22] (\new_sboxw[22] ), .\new_sboxw[23] (\new_sboxw[23] ), 
            .\enc_new_block[57] (enc_new_block[57]), .\round_logic.mixcolumns_block_39__N_1197[2] (\round_logic.mixcolumns_block_39__N_1197 [2]), 
            .\round_logic.mixcolumns_block_47__N_1397[6] (\round_logic.mixcolumns_block_47__N_1397 [6]), 
            .\round_logic.mixcolumns_block_15__N_1453[6] (\round_logic.mixcolumns_block_15__N_1453 [6]), 
            .\round_logic.mixcolumns_block_111__N_1285[5] (\round_logic.mixcolumns_block_111__N_1285 [5]), 
            .\round_logic.mixcolumns_block_79__N_1341[5] (\round_logic.mixcolumns_block_79__N_1341 [5]), 
            .n9638(n9638), .\enc_new_block[32] (enc_new_block[32]), .\round_logic.mixcolumns_block_7__N_1245[7] (\round_logic.mixcolumns_block_7__N_1245 [7]), 
            .\round_logic.mixcolumns_block_47__N_1397[5] (\round_logic.mixcolumns_block_47__N_1397 [5]), 
            .\round_logic.mixcolumns_block_15__N_1453[5] (\round_logic.mixcolumns_block_15__N_1453 [5]), 
            .\enc_new_block[43] (enc_new_block[43]), .\enc_new_block[11] (enc_new_block[11]), 
            .n9636(n9636), .\enc_new_block[107] (enc_new_block[107]), .\enc_new_block[75] (enc_new_block[75]), 
            .\enc_new_block[72] (enc_new_block[72]), .\round_logic.mixcolumns_block_15__N_1453[2] (\round_logic.mixcolumns_block_15__N_1453 [2]), 
            .\enc_new_block[42] (enc_new_block[42]), .\enc_new_block[10] (enc_new_block[10]), 
            .n9634(n9634), .\enc_new_block[106] (enc_new_block[106]), .\enc_new_block[74] (enc_new_block[74]), 
            .\round_logic.mixcolumns_block_111__N_1285[2] (\round_logic.mixcolumns_block_111__N_1285 [2]), 
            .\round_logic.mixcolumns_block_79__N_1341[2] (\round_logic.mixcolumns_block_79__N_1341 [2]), 
            .n9632(n9632), .\round_logic.mixcolumns_block_47__N_1397[2] (\round_logic.mixcolumns_block_47__N_1397 [2]), 
            .\round_key_gen.trw[2] (\round_key_gen.trw [2]), .\enc_new_block[26] (enc_new_block[26]), 
            .\enc_new_block[8] (enc_new_block[8]), .n9630(n9630), .\enc_new_block[104] (enc_new_block[104]), 
            .\enc_new_block[29] (enc_new_block[29]), .\round_logic.mixcolumns_block_7__N_1245[0] (\round_logic.mixcolumns_block_7__N_1245 [0]), 
            .\round_logic.mixcolumns_block_103__N_1101[0] (\round_logic.mixcolumns_block_103__N_1101 [0]), 
            .n9628(n9628), .\enc_new_block[31] (enc_new_block[31]), .\enc_new_block[64] (enc_new_block[64]), 
            .\round_logic.mixcolumns_block_39__N_1197[0] (\round_logic.mixcolumns_block_39__N_1197 [0]), 
            .\round_logic.mixcolumns_block_39__N_1197[7] (\round_logic.mixcolumns_block_39__N_1197 [7]), 
            .\round_logic.mixcolumns_block_103__N_1101[7] (\round_logic.mixcolumns_block_103__N_1101 [7]), 
            .n9626(n9626), .\round_logic.mixcolumns_block_71__N_1149[7] (\round_logic.mixcolumns_block_71__N_1149 [7]), 
            .\round_logic.mixcolumns_block_7__N_1245[6] (\round_logic.mixcolumns_block_7__N_1245 [6]), 
            .\round_logic.mixcolumns_block_103__N_1101[6] (\round_logic.mixcolumns_block_103__N_1101 [6]), 
            .n9624(n9624), .\round_logic.mixcolumns_block_71__N_1149[6] (\round_logic.mixcolumns_block_71__N_1149 [6]), 
            .\round_logic.mixcolumns_block_39__N_1197[6] (\round_logic.mixcolumns_block_39__N_1197 [6]), 
            .\round_logic.mixcolumns_block_7__N_1245[5] (\round_logic.mixcolumns_block_7__N_1245 [5]), 
            .\round_logic.mixcolumns_block_103__N_1101[5] (\round_logic.mixcolumns_block_103__N_1101 [5]), 
            .n9622(n9622), .\round_logic.mixcolumns_block_71__N_1149[5] (\round_logic.mixcolumns_block_71__N_1149 [5]), 
            .\round_logic.mixcolumns_block_39__N_1197[5] (\round_logic.mixcolumns_block_39__N_1197 [5]), 
            .\enc_new_block[35] (enc_new_block[35]), .\enc_new_block[3] (enc_new_block[3]), 
            .n9620(n9620), .\enc_new_block[99] (enc_new_block[99]), .\enc_new_block[34] (enc_new_block[34]), 
            .\enc_new_block[2] (enc_new_block[2]), .n9618(n9618), .\enc_new_block[98] (enc_new_block[98]), 
            .\enc_new_block[66] (enc_new_block[66]), .\round_logic.mixcolumns_block_7__N_1245[2] (\round_logic.mixcolumns_block_7__N_1245 [2]), 
            .\round_logic.mixcolumns_block_103__N_1101[2] (\round_logic.mixcolumns_block_103__N_1101 [2]), 
            .n9616(n9616), .\enc_new_block[63] (enc_new_block[63]), .\round_logic.mixcolumns_block_71__N_1149[2] (\round_logic.mixcolumns_block_71__N_1149 [2]), 
            .\enc_new_block[0] (enc_new_block[0]), .n8532(n8532), .\enc_new_block[96] (enc_new_block[96]), 
            .\enc_new_block[90] (enc_new_block[90]), .\enc_new_block[93] (enc_new_block[93]), 
            .\enc_new_block[94] (enc_new_block[94]), .\enc_new_block[95] (enc_new_block[95]), 
            .\enc_new_block[122] (enc_new_block[122]), .\enc_new_block[27] (enc_new_block[27]), 
            .\enc_new_block[28] (enc_new_block[28]), .\enc_new_block[30] (enc_new_block[30]), 
            .\block_reg[0][31] (\block_reg[0] [31]), .\enc_new_block[59] (enc_new_block[59]), 
            .\enc_new_block[60] (enc_new_block[60]), .\enc_new_block[61] (enc_new_block[61]), 
            .\enc_new_block[62] (enc_new_block[62]), .\block_reg[0][30] (\block_reg[0] [30]), 
            .\block_reg[0][28] (\block_reg[0] [28]), .\block_reg[0][26] (\block_reg[0] [26]), 
            .\enc_new_block[89] (enc_new_block[89]), .\enc_new_block[91] (enc_new_block[91]), 
            .\enc_new_block[92] (enc_new_block[92]), .block_w2_we_N_1489(n6364[2]), 
            .\block_reg[0][24] (\block_reg[0] [24]), .\round_key_gen.trw[0] (\round_key_gen.trw [0]), 
            .\block_reg[0][21] (\block_reg[0] [21]), .\enc_new_block[125] (enc_new_block[125]), 
            .\block_reg[0][16] (\block_reg[0] [16]), .\new_sboxw[16] (\new_sboxw[16] ), 
            .\block_reg[0][15] (\block_reg[0] [15]), .\enc_new_block[127] (enc_new_block[127]), 
            .\round_key_gen.trw[23] (\round_key_gen.trw [23]), .\block_reg[0][14] (\block_reg[0] [14]), 
            .\round_key_gen.trw[22] (\round_key_gen.trw [22]), .\block_reg[0][13] (\block_reg[0] [13]), 
            .\round_key_gen.trw[21] (\round_key_gen.trw [21]), .\block_reg[0][10] (\block_reg[0] [10]), 
            .\round_key_gen.trw[18] (\round_key_gen.trw [18]), .\block_reg[0][8] (\block_reg[0] [8]), 
            .\round_key_gen.trw[16] (\round_key_gen.trw [16]), .\block_reg[0][7] (\block_reg[0] [7]), 
            .n9676(n9676), .n9674(n9674), .\enc_new_block[126] (enc_new_block[126]), 
            .n9672(n9672), .n9670(n9670), .\enc_new_block[124] (enc_new_block[124]), 
            .n9668(n9668), .\enc_new_block[123] (enc_new_block[123]), .n9666(n9666), 
            .\enc_new_block[25] (enc_new_block[25]), .n9664(n9664), .\enc_new_block[121] (enc_new_block[121]), 
            .\block_new_127__N_1645[125] (block_new_127__N_1645[125]), .\block_new_127__N_1645[123] (block_new_127__N_1645[123]), 
            .\block_new_127__N_1645[121] (block_new_127__N_1645[121]), .\block_new_127__N_1645[119] (block_new_127__N_1645[119]), 
            .\block_reg[1][24] (\block_reg[1] [24]), .\block_new_127__N_1645[118] (block_new_127__N_1645[118]), 
            .\block_new_127__N_1645[116] (block_new_127__N_1645[116]), .\block_new_127__N_1645[115] (block_new_127__N_1645[115]), 
            .\block_new_127__N_1645[114] (block_new_127__N_1645[114]), .\block_new_127__N_1645[113] (block_new_127__N_1645[113]), 
            .\block_new_127__N_1645[108] (block_new_127__N_1645[108]), .\block_reg[1][16] (\block_reg[1] [16]), 
            .\block_reg[1][15] (\block_reg[1] [15]), .n33848(n33848), .\block_reg[1][14] (\block_reg[1] [14]), 
            .\block_reg[1][13] (\block_reg[1] [13]), .\block_new_127__N_1645[107] (block_new_127__N_1645[107]), 
            .\block_new_127__N_1645[105] (block_new_127__N_1645[105]), .\block_new_127__N_1645[102] (block_new_127__N_1645[102]), 
            .\block_reg[1][10] (\block_reg[1] [10]), .\block_new_127__N_1645[99] (block_new_127__N_1645[99]), 
            .\block_new_127__N_1645[98] (block_new_127__N_1645[98]), .\block_new_127__N_1645[97] (block_new_127__N_1645[97]), 
            .\block_reg[1][8] (\block_reg[1] [8]), .\block_reg[2][3] (\block_reg[2] [3]), 
            .enc_round_nr({enc_round_nr}), .\block_new_127__N_1645[92] (block_new_127__N_1645[92]), 
            .\block_new_127__N_1645[91] (block_new_127__N_1645[91]), .\block_new_127__N_1645[89] (block_new_127__N_1645[89]), 
            .\block_new_127__N_1645[87] (block_new_127__N_1645[87]), .\block_new_127__N_1645[86] (block_new_127__N_1645[86]), 
            .\block_new_127__N_1645[85] (block_new_127__N_1645[85]), .\block_new_127__N_1645[84] (block_new_127__N_1645[84]), 
            .\block_reg[1][2] (\block_reg[1] [2]), .\block_new_127__N_1645[83] (block_new_127__N_1645[83]), 
            .\block_new_127__N_1645[82] (block_new_127__N_1645[82]), .\block_new_127__N_1645[81] (block_new_127__N_1645[81]), 
            .\block_new_127__N_1645[76] (block_new_127__N_1645[76]), .\block_reg[2][31] (\block_reg[2] [31]), 
            .\block_new_127__N_1645[75] (block_new_127__N_1645[75]), .\block_new_127__N_1645[73] (block_new_127__N_1645[73]), 
            .\block_new_127__N_1645[71] (block_new_127__N_1645[71]), .\block_new_127__N_1645[70] (block_new_127__N_1645[70]), 
            .\block_reg[2][26] (\block_reg[2] [26]), .n33913(n33913), .n28773(n28773), 
            .\block_reg[2][24] (\block_reg[2] [24]), .\block_reg[2][23] (\block_reg[2] [23]), 
            .\block_new_127__N_1645[69] (block_new_127__N_1645[69]), .\block_reg[2][22] (\block_reg[2] [22]), 
            .\block_reg[2][21] (\block_reg[2] [21]), .\block_reg[2][20] (\block_reg[2] [20]), 
            .\block_reg[2][16] (\block_reg[2] [16]), .\block_reg[2][15] (\block_reg[2] [15]), 
            .\block_reg[2][14] (\block_reg[2] [14]), .\block_new_127__N_1645[68] (block_new_127__N_1645[68]), 
            .\block_new_127__N_1645[67] (block_new_127__N_1645[67]), .\block_reg[2][13] (\block_reg[2] [13]), 
            .\block_new_127__N_1645[65] (block_new_127__N_1645[65]), .\block_reg[2][10] (\block_reg[2] [10]), 
            .\block_new_127__N_1645[64] (block_new_127__N_1645[64]), .\block_reg[2][8] (\block_reg[2] [8]), 
            .\block_reg[2][6] (\block_reg[2] [6]), .n5(n5), .round_ctr_we(round_ctr_we), 
            .n33915(n33915), .\block_new_127__N_1645[62] (block_new_127__N_1645[62]), 
            .\block_new_127__N_1645[61] (block_new_127__N_1645[61]), .\key_mem_ctrl.num_rounds[2] (\key_mem_ctrl.num_rounds[2] ), 
            .n4(n4), .\block_new_127__N_1645[12] (block_new_127__N_1645[12]), 
            .\block_new_127__N_1645[60] (block_new_127__N_1645[60]), .\block_new_127__N_1645[10] (block_new_127__N_1645[10]), 
            .\block_new_127__N_1645[7] (block_new_127__N_1645[7]), .\block_new_127__N_1645[59] (block_new_127__N_1645[59]), 
            .\block_new_127__N_1645[5] (block_new_127__N_1645[5]), .\block_new_127__N_1645[4] (block_new_127__N_1645[4]), 
            .\block_new_127__N_1645[57] (block_new_127__N_1645[57]), .\block_reg[2][0] (\block_reg[2] [0]), 
            .\block_reg[3][31] (\block_reg[3] [31]), .\block_reg[3][29] (\block_reg[3] [29]), 
            .\block_new_127__N_1645[3] (block_new_127__N_1645[3]), .\block_new_127__N_1645[2] (block_new_127__N_1645[2]), 
            .\block_reg[3][26] (\block_reg[3] [26]), .\block_new_127__N_1645[1] (block_new_127__N_1645[1]), 
            .\block_reg[3][24] (\block_reg[3] [24]), .\block_reg[3][23] (\block_reg[3] [23]), 
            .\block_new_127__N_1645[51] (block_new_127__N_1645[51]), .\block_reg[3][22] (\block_reg[3] [22]), 
            .\block_new_127__N_1645[50] (block_new_127__N_1645[50]), .\block_new_127__N_1645[49] (block_new_127__N_1645[49]), 
            .\block_reg[3][18] (\block_reg[3] [18]), .\block_new_127__N_1645[44] (block_new_127__N_1645[44]), 
            .\block_new_127__N_1645[43] (block_new_127__N_1645[43]), .\block_new_127__N_1645[41] (block_new_127__N_1645[41]), 
            .\block_reg[3][16] (\block_reg[3] [16]), .\block_reg[3][15] (\block_reg[3] [15]), 
            .\block_new_127__N_1645[39] (block_new_127__N_1645[39]), .\block_new_127__N_1645[37] (block_new_127__N_1645[37]), 
            .\block_new_127__N_1645[36] (block_new_127__N_1645[36]), .\block_new_127__N_1645[34] (block_new_127__N_1645[34]), 
            .\block_reg[3][13] (\block_reg[3] [13]), .\block_new_127__N_1645[33] (block_new_127__N_1645[33]), 
            .\block_new_127__N_1645[30] (block_new_127__N_1645[30]), .\block_reg[3][11] (\block_reg[3] [11]), 
            .\block_new_127__N_1645[28] (block_new_127__N_1645[28]), .\block_new_127__N_1645[27] (block_new_127__N_1645[27]), 
            .\block_reg[3][9] (\block_reg[3] [9]), .\block_new_127__N_1645[25] (block_new_127__N_1645[25]), 
            .\block_reg[3][8] (\block_reg[3] [8]), .\block_reg[3][6] (\block_reg[3] [6]), 
            .\block_new_127__N_1645[21] (block_new_127__N_1645[21]), .\block_new_127__N_1645[20] (block_new_127__N_1645[20]), 
            .\block_new_127__N_1645[19] (block_new_127__N_1645[19]), .\block_new_127__N_1645[17] (block_new_127__N_1645[17]), 
            .\block_new_127__N_1645[14] (block_new_127__N_1645[14]), .\block_reg[3][0] (\block_reg[3] [0])) /* synthesis syn_module_defined=1 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(116[22] 132[32])
    aes_decipher_block dec_block (.dec_new_block({dec_new_block}), .round_key({round_key}), 
            .clk_c(clk_c), .tmp_sboxw({tmp_sboxw}), .dec_round_nr({Open_3, 
            Open_4, Open_5, \dec_round_nr[0] }), .round_ctr_we(round_ctr_we_adj_128), 
            .round_ctr_new({Open_6, Open_7, Open_8, \round_ctr_new[0] }), 
            .n6347({enc_ctrl_new_2__N_1045, n6347[2:0]}), .encdec_reg(encdec_reg), 
            .\aes_core_ctrl_new_1__N_858[1] (\aes_core_ctrl_new_1__N_858[1] ), 
            .n28773(n28773), .\enc_round_nr[3] (enc_round_nr[3]), .block_w3_we_N_1490(n6364[3]), 
            .n4(n4), .n33858(n33858), .n149(n149), .block_new_127__N_1645({Open_9, 
            Open_10, Open_11, Open_12, Open_13, Open_14, Open_15, 
            Open_16, Open_17, Open_18, Open_19, Open_20, Open_21, 
            Open_22, Open_23, Open_24, Open_25, Open_26, Open_27, 
            Open_28, Open_29, Open_30, Open_31, Open_32, Open_33, 
            Open_34, Open_35, Open_36, Open_37, Open_38, Open_39, 
            Open_40, Open_41, Open_42, Open_43, Open_44, Open_45, 
            Open_46, Open_47, Open_48, Open_49, Open_50, Open_51, 
            Open_52, Open_53, Open_54, Open_55, Open_56, Open_57, 
            Open_58, Open_59, Open_60, Open_61, Open_62, Open_63, 
            Open_64, Open_65, Open_66, Open_67, Open_68, Open_69, 
            Open_70, Open_71, Open_72, Open_73, Open_74, Open_75, 
            Open_76, Open_77, Open_78, Open_79, Open_80, Open_81, 
            Open_82, Open_83, Open_84, Open_85, Open_86, Open_87, 
            Open_88, Open_89, Open_90, Open_91, Open_92, Open_93, 
            Open_94, Open_95, Open_96, block_new_127__N_1645[39], Open_97, 
            Open_98, Open_99, Open_100, Open_101, Open_102, Open_103, 
            Open_104, Open_105, Open_106, Open_107, Open_108, Open_109, 
            Open_110, Open_111, Open_112, Open_113, Open_114, Open_115, 
            Open_116, Open_117, Open_118, Open_119, Open_120, Open_121, 
            Open_122, Open_123, Open_124, Open_125, Open_126, Open_127, 
            Open_128, Open_129, Open_130, Open_131, Open_132, Open_133, 
            Open_134, Open_135}), .\block_new_127__N_1645[37] (block_new_127__N_1645[37]), 
            .\block_new_127__N_1645[36] (block_new_127__N_1645[36]), .\block_new_127__N_1645[34] (block_new_127__N_1645[34]), 
            .\block_new_127__N_1645[33] (block_new_127__N_1645[33]), .\block_new_127__N_1645[62] (block_new_127__N_1645[62]), 
            .\block_new_127__N_1645[61] (block_new_127__N_1645[61]), .\block_new_127__N_1645[60] (block_new_127__N_1645[60]), 
            .\block_new_127__N_1645[59] (block_new_127__N_1645[59]), .\block_new_127__N_1645[57] (block_new_127__N_1645[57]), 
            .\block_new_127__N_1645[87] (block_new_127__N_1645[87]), .\block_new_127__N_1645[86] (block_new_127__N_1645[86]), 
            .\block_new_127__N_1645[85] (block_new_127__N_1645[85]), .\block_new_127__N_1645[84] (block_new_127__N_1645[84]), 
            .\block_new_127__N_1645[83] (block_new_127__N_1645[83]), .\block_new_127__N_1645[82] (block_new_127__N_1645[82]), 
            .\block_new_127__N_1645[81] (block_new_127__N_1645[81]), .\block_new_127__N_1645[108] (block_new_127__N_1645[108]), 
            .\block_new_127__N_1645[107] (block_new_127__N_1645[107]), .\block_new_127__N_1645[105] (block_new_127__N_1645[105]), 
            .\block_new_127__N_1645[7] (block_new_127__N_1645[7]), .\block_new_127__N_1645[5] (block_new_127__N_1645[5]), 
            .\block_new_127__N_1645[4] (block_new_127__N_1645[4]), .\block_new_127__N_1645[3] (block_new_127__N_1645[3]), 
            .\block_new_127__N_1645[2] (block_new_127__N_1645[2]), .\enc_round_nr[1] (enc_round_nr[1]), 
            .\muxed_round_nr[1] (muxed_round_nr[1]), .\block_new_127__N_1645[1] (block_new_127__N_1645[1]), 
            .\block_new_127__N_1645[30] (block_new_127__N_1645[30]), .new_sboxw({new_sboxw}), 
            .\block_new_127__N_1645[28] (block_new_127__N_1645[28]), .\block_new_127__N_1645[27] (block_new_127__N_1645[27]), 
            .\block_new_127__N_1645[25] (block_new_127__N_1645[25]), .\block_reg[0] ({\block_reg[0] }), 
            .\block_new_127__N_1645[51] (block_new_127__N_1645[51]), .\block_new_127__N_1645[50] (block_new_127__N_1645[50]), 
            .\block_new_127__N_1645[49] (block_new_127__N_1645[49]), .dec_ready(dec_ready), 
            .dec_ctrl_we(dec_ctrl_we), .\block_new_127__N_1645[76] (block_new_127__N_1645[76]), 
            .\block_new_127__N_1645[125] (block_new_127__N_1645[125]), .\block_new_127__N_1645[123] (block_new_127__N_1645[123]), 
            .\key_mem_ctrl.num_rounds[2] (\key_mem_ctrl.num_rounds[2] ), .\muxed_round_nr[3] (muxed_round_nr[3]), 
            .\enc_round_nr[2] (enc_round_nr[2]), .\muxed_round_nr[2] (muxed_round_nr[2]), 
            .\block_new_127__N_1645[121] (block_new_127__N_1645[121]), .\block_new_127__N_1645[21] (block_new_127__N_1645[21]), 
            .\block_new_127__N_1645[20] (block_new_127__N_1645[20]), .\block_new_127__N_1645[19] (block_new_127__N_1645[19]), 
            .\block_new_127__N_1645[17] (block_new_127__N_1645[17]), .\block_new_127__N_1645[44] (block_new_127__N_1645[44]), 
            .\block_new_127__N_1645[43] (block_new_127__N_1645[43]), .\block_new_127__N_1645[41] (block_new_127__N_1645[41]), 
            .\block_new_127__N_1645[71] (block_new_127__N_1645[71]), .\block_new_127__N_1645[70] (block_new_127__N_1645[70]), 
            .\block_new_127__N_1645[69] (block_new_127__N_1645[69]), .\block_new_127__N_1645[68] (block_new_127__N_1645[68]), 
            .\block_new_127__N_1645[67] (block_new_127__N_1645[67]), .\block_new_127__N_1645[65] (block_new_127__N_1645[65]), 
            .\block_new_127__N_1645[64] (block_new_127__N_1645[64]), .\block_new_127__N_1645[92] (block_new_127__N_1645[92]), 
            .\block_new_127__N_1645[91] (block_new_127__N_1645[91]), .\block_new_127__N_1645[89] (block_new_127__N_1645[89]), 
            .\block_new_127__N_1645[119] (block_new_127__N_1645[119]), .\block_new_127__N_1645[118] (block_new_127__N_1645[118]), 
            .\block_new_127__N_1645[116] (block_new_127__N_1645[116]), .\block_new_127__N_1645[115] (block_new_127__N_1645[115]), 
            .\block_new_127__N_1645[114] (block_new_127__N_1645[114]), .\block_new_127__N_1645[113] (block_new_127__N_1645[113]), 
            .\block_new_127__N_1645[14] (block_new_127__N_1645[14]), .\block_new_127__N_1645[12] (block_new_127__N_1645[12]), 
            .\block_new_127__N_1645[10] (block_new_127__N_1645[10]), .\block_new_127__N_1645[75] (block_new_127__N_1645[75]), 
            .\block_new_127__N_1645[73] (block_new_127__N_1645[73]), .\block_new_127__N_1645[102] (block_new_127__N_1645[102]), 
            .\block_new_127__N_1645[99] (block_new_127__N_1645[99]), .\block_new_127__N_1645[98] (block_new_127__N_1645[98]), 
            .\block_new_127__N_1645[97] (block_new_127__N_1645[97]), .n14934(n14934), 
            .dec_ctrl_new_2__N_2032(dec_ctrl_new_2__N_2032), .n33848(n33848), 
            .n33846(n33846), .\block_reg[1] ({\block_reg[1] }), .\block_reg[3] ({\block_reg[3] }), 
            .\round_ctr_new[3] (\round_ctr_new[3] ), .n33942(n33942), .n33913(n33913), 
            .enc_ready(enc_ready), .n6428(n6428), .\block_reg[2] ({\block_reg[2] }), 
            .n14930(n14930), .n33909(n33909), .n14939(n14939), .n152(n152)) /* synthesis syn_module_defined=1 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(135[22] 148[32])
    
endmodule
//
// Verilog Description of module aes_key_mem
//

module aes_key_mem (n33952, \muxed_round_nr[1] , \round_key_gen.trw[2] , 
            n33860, \key_reg[0] , n11, \round_key_gen.trw[1] , n35835, 
            clk_c, GND_net, \round_key_gen.trw[0] , \new_sboxw[23] , 
            \new_sboxw[22] , \key_mem_ctrl.num_rounds[2] , \key_reg[3] , 
            \key_reg[2] , \key_reg[1] , n11_adj_1, \new_sboxw[21] , 
            \key_reg[5] , \new_sboxw[20] , \new_sboxw[19] , n11_adj_2, 
            n11_adj_3, n15316, \key_reg[6] , \round_key_gen.trw[8] , 
            n15429, \round_key_gen.trw[9] , n15489, \round_key_gen.trw[10] , 
            n15549, \round_key_gen.trw[3] , \round_key_gen.trw[11] , n15609, 
            n11_adj_4, \round_key_gen.trw[4] , \round_key_gen.trw[12] , 
            n15669, \round_key_gen.trw[5] , \round_key_gen.trw[13] , n15729, 
            \round_key_gen.trw[6] , \round_key_gen.trw[14] , n15789, \round_key_gen.trw[7] , 
            \round_key_gen.trw[15] , n15849, \round_key_gen.trw[16] , 
            n11_adj_5, n15909, n11_adj_6, \round_key_gen.trw[17] , n15969, 
            \round_key_gen.trw[18] , n16029, \new_sboxw[18] , \round_key_gen.trw[19] , 
            \new_sboxw[17] , n11_adj_7, n16089, \round_key_gen.trw[20] , 
            n16149, \round_key_gen.trw[21] , n11_adj_8, n16209, \round_key_gen.trw[22] , 
            n16269, \round_key_gen.trw[23] , n16329, \new_sboxw[16] , 
            n11_adj_9, n16389, n11_adj_10, n16449, n11_adj_11, n16509, 
            n16569, n11_adj_12, n11_adj_13, n16629, n16689, n11_adj_14, 
            n16749, n16809, n11_adj_15, n16869, n11_adj_16, n16929, 
            n11_adj_17, n16989, n17049, n17109, n17169, n11_adj_18, 
            n17229, n11_adj_19, n11_adj_20, \key_reg[4] , n11_adj_21, 
            n11_adj_22, n11_adj_23, n11_adj_24, n11_adj_25, n11_adj_26, 
            n11_adj_27, n11_adj_28, n11_adj_29, n11_adj_30, n11_adj_31, 
            n11_adj_32, n11_adj_33, \key_mem[14] , n11_adj_34, n5, 
            init_state, n11_adj_35, n11_adj_36, n11_adj_37, n11_adj_38, 
            n11_adj_39, n11_adj_40, n11_adj_41, \muxed_sboxw[16] , \muxed_sboxw[17] , 
            \muxed_sboxw[18] , \muxed_sboxw[19] , \muxed_sboxw[20] , n11_adj_42, 
            \muxed_sboxw[21] , \muxed_sboxw[22] , \muxed_sboxw[23] , key_ready, 
            n11_adj_43, n11_adj_44, n11_adj_45, n11_adj_46, reset_n_c, 
            n11_adj_47, n11_adj_48, n11_adj_49, n11_adj_50, n11_adj_51, 
            n11_adj_52, n11_adj_53, n11_adj_54, n11_adj_55, n11_adj_56, 
            n11_adj_57, n11_adj_58, n11_adj_59, n11_adj_60, n11_adj_61, 
            n11_adj_62, n11_adj_63, n11_adj_64, n11_adj_65, n11_adj_66, 
            n11_adj_67, n11_adj_68, n11_adj_69, n11_adj_70, n11_adj_71, 
            n11_adj_72, n11_adj_73, n11_adj_74, n11_adj_75, n11_adj_76, 
            n11_adj_77, \muxed_round_nr[3] , round_key, n11_adj_78, 
            n11_adj_79, n11_adj_80, n11_adj_81, n11_adj_82, n11_adj_83, 
            n11_adj_84, n11_adj_85, n11_adj_86, n11_adj_87, n11_adj_88, 
            n11_adj_89, \key_reg[7] , n11_adj_90, n11_adj_91, n11_adj_92, 
            n11_adj_93, n11_adj_94, n11_adj_95, \muxed_round_nr[2] , 
            n33343, n33344, n33345, n33346, n33347, n33348, n33349, 
            n33351, n33352, n33353, n33354, n33356, n33357, n33358, 
            n33359, n33360, n33362, n33363, n33364, n33365, n11_adj_96, 
            n33366, n33368, n33369, n33370, n33371, n11_adj_97, 
            n33372, n33373, n33375, n33376, n33378, n33381, n33383, 
            n33385, n33388, n33390, n11_adj_98, n11_adj_99, n11_adj_100, 
            n33392, n11_adj_101, n17224, n17164, n17104, n11_adj_102, 
            n17044, n16984, n16924, n16864, n16804, n16744, n16684, 
            n16624, n11_adj_103, n16564, n16504, n16444, n16384, 
            n16324, n16264, n16204, n16144, n16084, n11_adj_104, 
            n16024, n15964, n15904, n15844, n15784, n15724, n15664, 
            n15604, n15544, n15484, n15424, n11_adj_105, n11_adj_106, 
            n11_adj_107, n11_adj_108, n11_adj_109, n11_adj_110, n11_adj_111, 
            n33394, n11_adj_112, n33396, n33397, n33399, n33401, 
            n11_adj_113, n33403, n11_adj_114, maxfan_replicated_net_23, 
            n11_adj_115, n33404, n33407, n33408, n33410, n11_adj_116, 
            n33412, n33414, n33415, n33416, n11_adj_117, n33417, 
            n33418, n33419, n33420, n33421, n33422, n33423, n33424, 
            n33425, n33426, n33427, n33428, n33429, n33430, n11_adj_118, 
            n11_adj_119, n11_adj_120, n11_adj_121, n11_adj_122, \prev_key1_new_127__N_4787[1] , 
            \prev_key1_new_127__N_4787[2] , \prev_key1_new_127__N_4787[3] , 
            \prev_key1_new_127__N_4787[4] , \prev_key1_new_127__N_4787[5] , 
            \prev_key1_new_127__N_4787[6] , \prev_key1_new_127__N_4787[7] , 
            \prev_key1_new_127__N_4787[8] , \prev_key1_new_127__N_4787[9] , 
            \prev_key1_new_127__N_4787[10] , \prev_key1_new_127__N_4787[11] , 
            \prev_key1_new_127__N_4787[12] , \prev_key1_new_127__N_4787[13] , 
            \prev_key1_new_127__N_4787[14] , \prev_key1_new_127__N_4787[15] , 
            \prev_key1_new_127__N_4787[16] , \prev_key1_new_127__N_4787[17] , 
            \prev_key1_new_127__N_4787[18] , \prev_key1_new_127__N_4787[19] , 
            \prev_key1_new_127__N_4787[20] , \prev_key1_new_127__N_4787[21] , 
            \prev_key1_new_127__N_4787[22] , \prev_key1_new_127__N_4787[23] , 
            \prev_key1_new_127__N_4787[24] , \prev_key1_new_127__N_4787[25] , 
            \prev_key1_new_127__N_4787[26] , \prev_key1_new_127__N_4787[27] , 
            \prev_key1_new_127__N_4787[28] , \prev_key1_new_127__N_4787[29] , 
            \prev_key1_new_127__N_4787[30] , \prev_key1_new_127__N_4787[31] , 
            \prev_key1_new_127__N_4787[32] , \prev_key1_new_127__N_4787[33] , 
            \prev_key1_new_127__N_4787[34] , \prev_key1_new_127__N_4787[35] , 
            \prev_key1_new_127__N_4787[36] , \prev_key1_new_127__N_4787[37] , 
            \prev_key1_new_127__N_4787[38] , \prev_key1_new_127__N_4787[39] , 
            \prev_key1_new_127__N_4787[40] , \prev_key1_new_127__N_4787[41] , 
            \prev_key1_new_127__N_4787[42] , \prev_key1_new_127__N_4787[43] , 
            \prev_key1_new_127__N_4787[44] , \prev_key1_new_127__N_4787[45] , 
            \prev_key1_new_127__N_4787[46] , \prev_key1_new_127__N_4787[47] , 
            \prev_key1_new_127__N_4787[48] , \prev_key1_new_127__N_4787[49] , 
            \prev_key1_new_127__N_4787[50] , \prev_key1_new_127__N_4787[51] , 
            \prev_key1_new_127__N_4787[52] , \prev_key1_new_127__N_4787[53] , 
            \prev_key1_new_127__N_4787[54] , \prev_key1_new_127__N_4787[55] , 
            \prev_key1_new_127__N_4787[56] , \prev_key1_new_127__N_4787[57] , 
            \prev_key1_new_127__N_4787[58] , \prev_key1_new_127__N_4787[59] , 
            \prev_key1_new_127__N_4787[60] , \prev_key1_new_127__N_4787[61] , 
            \prev_key1_new_127__N_4787[62] , \prev_key1_new_127__N_4787[63] , 
            n33431, n33432, n11_adj_123, n33433, n33434, n33436, 
            n33441, n33446, n33448, n33449, n33450, n33451, n33452, 
            n33453, n33454, n33455, n33456, n33457, n33458, n33459, 
            n33460, n33461, n11_adj_124, n33462, n33463, n33336, 
            n33435, n33437, n33438, n33439, n33440, n33442, n33443, 
            n33444, n33445, n33447, n33337, n33338, n33339, n33340, 
            n33341, n33342, n33350, n33355, n33361, n33367, n33374, 
            n33377, n33379, n33380, n33382, n33384, n33386, n11_adj_125, 
            n33387, n33389, n33391, n33393, n33395, n33398, n33400, 
            n33402, n33405, n33406, n33409, n33411, n33413, n11_adj_126, 
            n2531, n8532, n9616, n9618, n9620, n9622, n9624, n9626, 
            n9628, n9630, n9632, n9634, n9636, n9638, n9640, n9642, 
            n9644, n9646, n9648, n9650, n9652, n9654, n9656, n9658, 
            n9660, n9662, n11_adj_127, n9664, n9666, n9668, n9670, 
            n9672, n9674, n9676, \key_mem_ctrl_new_2__N_4928[0] , block_w3_we_N_1490, 
            block_w2_we_N_1489) /* synthesis syn_module_defined=1 */ ;
    input n33952;
    input \muxed_round_nr[1] ;
    output \round_key_gen.trw[2] ;
    output n33860;
    input [31:0]\key_reg[0] ;
    output n11;
    output \round_key_gen.trw[1] ;
    input n35835;
    input clk_c;
    input GND_net;
    output \round_key_gen.trw[0] ;
    input \new_sboxw[23] ;
    input \new_sboxw[22] ;
    input \key_mem_ctrl.num_rounds[2] ;
    input [31:0]\key_reg[3] ;
    input [31:0]\key_reg[2] ;
    input [31:0]\key_reg[1] ;
    output n11_adj_1;
    input \new_sboxw[21] ;
    input [31:0]\key_reg[5] ;
    input \new_sboxw[20] ;
    input \new_sboxw[19] ;
    output n11_adj_2;
    output n11_adj_3;
    output n15316;
    input [31:0]\key_reg[6] ;
    output \round_key_gen.trw[8] ;
    output n15429;
    output \round_key_gen.trw[9] ;
    output n15489;
    output \round_key_gen.trw[10] ;
    output n15549;
    output \round_key_gen.trw[3] ;
    output \round_key_gen.trw[11] ;
    output n15609;
    output n11_adj_4;
    output \round_key_gen.trw[4] ;
    output \round_key_gen.trw[12] ;
    output n15669;
    output \round_key_gen.trw[5] ;
    output \round_key_gen.trw[13] ;
    output n15729;
    output \round_key_gen.trw[6] ;
    output \round_key_gen.trw[14] ;
    output n15789;
    output \round_key_gen.trw[7] ;
    output \round_key_gen.trw[15] ;
    output n15849;
    output \round_key_gen.trw[16] ;
    output n11_adj_5;
    output n15909;
    output n11_adj_6;
    output \round_key_gen.trw[17] ;
    output n15969;
    output \round_key_gen.trw[18] ;
    output n16029;
    input \new_sboxw[18] ;
    output \round_key_gen.trw[19] ;
    input \new_sboxw[17] ;
    output n11_adj_7;
    output n16089;
    output \round_key_gen.trw[20] ;
    output n16149;
    output \round_key_gen.trw[21] ;
    output n11_adj_8;
    output n16209;
    output \round_key_gen.trw[22] ;
    output n16269;
    output \round_key_gen.trw[23] ;
    output n16329;
    input \new_sboxw[16] ;
    output n11_adj_9;
    output n16389;
    output n11_adj_10;
    output n16449;
    output n11_adj_11;
    output n16509;
    output n16569;
    output n11_adj_12;
    output n11_adj_13;
    output n16629;
    output n16689;
    output n11_adj_14;
    output n16749;
    output n16809;
    output n11_adj_15;
    output n16869;
    output n11_adj_16;
    output n16929;
    output n11_adj_17;
    output n16989;
    output n17049;
    output n17109;
    output n17169;
    output n11_adj_18;
    output n17229;
    output n11_adj_19;
    output n11_adj_20;
    input [31:0]\key_reg[4] ;
    output n11_adj_21;
    output n11_adj_22;
    output n11_adj_23;
    output n11_adj_24;
    output n11_adj_25;
    output n11_adj_26;
    output n11_adj_27;
    output n11_adj_28;
    output n11_adj_29;
    output n11_adj_30;
    output n11_adj_31;
    output n11_adj_32;
    output n11_adj_33;
    output [127:0]\key_mem[14] ;
    output n11_adj_34;
    input n5;
    input init_state;
    output n11_adj_35;
    output n11_adj_36;
    output n11_adj_37;
    output n11_adj_38;
    output n11_adj_39;
    output n11_adj_40;
    output n11_adj_41;
    output \muxed_sboxw[16] ;
    output \muxed_sboxw[17] ;
    output \muxed_sboxw[18] ;
    output \muxed_sboxw[19] ;
    output \muxed_sboxw[20] ;
    output n11_adj_42;
    output \muxed_sboxw[21] ;
    output \muxed_sboxw[22] ;
    output \muxed_sboxw[23] ;
    output key_ready;
    output n11_adj_43;
    output n11_adj_44;
    output n11_adj_45;
    output n11_adj_46;
    input reset_n_c;
    output n11_adj_47;
    output n11_adj_48;
    output n11_adj_49;
    output n11_adj_50;
    output n11_adj_51;
    output n11_adj_52;
    output n11_adj_53;
    output n11_adj_54;
    output n11_adj_55;
    output n11_adj_56;
    output n11_adj_57;
    output n11_adj_58;
    output n11_adj_59;
    output n11_adj_60;
    output n11_adj_61;
    output n11_adj_62;
    output n11_adj_63;
    output n11_adj_64;
    output n11_adj_65;
    output n11_adj_66;
    output n11_adj_67;
    output n11_adj_68;
    output n11_adj_69;
    output n11_adj_70;
    output n11_adj_71;
    output n11_adj_72;
    output n11_adj_73;
    output n11_adj_74;
    output n11_adj_75;
    output n11_adj_76;
    output n11_adj_77;
    input \muxed_round_nr[3] ;
    output [127:0]round_key;
    output n11_adj_78;
    output n11_adj_79;
    output n11_adj_80;
    output n11_adj_81;
    output n11_adj_82;
    output n11_adj_83;
    output n11_adj_84;
    output n11_adj_85;
    output n11_adj_86;
    output n11_adj_87;
    output n11_adj_88;
    output n11_adj_89;
    input [31:0]\key_reg[7] ;
    output n11_adj_90;
    output n11_adj_91;
    output n11_adj_92;
    output n11_adj_93;
    output n11_adj_94;
    output n11_adj_95;
    input \muxed_round_nr[2] ;
    input n33343;
    input n33344;
    input n33345;
    input n33346;
    input n33347;
    input n33348;
    input n33349;
    input n33351;
    input n33352;
    input n33353;
    input n33354;
    input n33356;
    input n33357;
    input n33358;
    input n33359;
    input n33360;
    input n33362;
    input n33363;
    input n33364;
    input n33365;
    output n11_adj_96;
    input n33366;
    input n33368;
    input n33369;
    input n33370;
    input n33371;
    output n11_adj_97;
    input n33372;
    input n33373;
    input n33375;
    input n33376;
    input n33378;
    input n33381;
    input n33383;
    input n33385;
    input n33388;
    input n33390;
    output n11_adj_98;
    output n11_adj_99;
    output n11_adj_100;
    input n33392;
    output n11_adj_101;
    output n17224;
    output n17164;
    output n17104;
    output n11_adj_102;
    output n17044;
    output n16984;
    output n16924;
    output n16864;
    output n16804;
    output n16744;
    output n16684;
    output n16624;
    output n11_adj_103;
    output n16564;
    output n16504;
    output n16444;
    output n16384;
    output n16324;
    output n16264;
    output n16204;
    output n16144;
    output n16084;
    output n11_adj_104;
    output n16024;
    output n15964;
    output n15904;
    output n15844;
    output n15784;
    output n15724;
    output n15664;
    output n15604;
    output n15544;
    output n15484;
    output n15424;
    output n11_adj_105;
    output n11_adj_106;
    output n11_adj_107;
    output n11_adj_108;
    output n11_adj_109;
    output n11_adj_110;
    output n11_adj_111;
    input n33394;
    output n11_adj_112;
    input n33396;
    input n33397;
    input n33399;
    input n33401;
    output n11_adj_113;
    input n33403;
    output n11_adj_114;
    input maxfan_replicated_net_23;
    output n11_adj_115;
    input n33404;
    input n33407;
    input n33408;
    input n33410;
    output n11_adj_116;
    input n33412;
    input n33414;
    input n33415;
    input n33416;
    output n11_adj_117;
    input n33417;
    input n33418;
    input n33419;
    input n33420;
    input n33421;
    input n33422;
    input n33423;
    input n33424;
    input n33425;
    input n33426;
    input n33427;
    input n33428;
    input n33429;
    input n33430;
    output n11_adj_118;
    output n11_adj_119;
    output n11_adj_120;
    output n11_adj_121;
    output n11_adj_122;
    input \prev_key1_new_127__N_4787[1] ;
    input \prev_key1_new_127__N_4787[2] ;
    input \prev_key1_new_127__N_4787[3] ;
    input \prev_key1_new_127__N_4787[4] ;
    input \prev_key1_new_127__N_4787[5] ;
    input \prev_key1_new_127__N_4787[6] ;
    input \prev_key1_new_127__N_4787[7] ;
    input \prev_key1_new_127__N_4787[8] ;
    input \prev_key1_new_127__N_4787[9] ;
    input \prev_key1_new_127__N_4787[10] ;
    input \prev_key1_new_127__N_4787[11] ;
    input \prev_key1_new_127__N_4787[12] ;
    input \prev_key1_new_127__N_4787[13] ;
    input \prev_key1_new_127__N_4787[14] ;
    input \prev_key1_new_127__N_4787[15] ;
    input \prev_key1_new_127__N_4787[16] ;
    input \prev_key1_new_127__N_4787[17] ;
    input \prev_key1_new_127__N_4787[18] ;
    input \prev_key1_new_127__N_4787[19] ;
    input \prev_key1_new_127__N_4787[20] ;
    input \prev_key1_new_127__N_4787[21] ;
    input \prev_key1_new_127__N_4787[22] ;
    input \prev_key1_new_127__N_4787[23] ;
    input \prev_key1_new_127__N_4787[24] ;
    input \prev_key1_new_127__N_4787[25] ;
    input \prev_key1_new_127__N_4787[26] ;
    input \prev_key1_new_127__N_4787[27] ;
    input \prev_key1_new_127__N_4787[28] ;
    input \prev_key1_new_127__N_4787[29] ;
    input \prev_key1_new_127__N_4787[30] ;
    input \prev_key1_new_127__N_4787[31] ;
    input \prev_key1_new_127__N_4787[32] ;
    input \prev_key1_new_127__N_4787[33] ;
    input \prev_key1_new_127__N_4787[34] ;
    input \prev_key1_new_127__N_4787[35] ;
    input \prev_key1_new_127__N_4787[36] ;
    input \prev_key1_new_127__N_4787[37] ;
    input \prev_key1_new_127__N_4787[38] ;
    input \prev_key1_new_127__N_4787[39] ;
    input \prev_key1_new_127__N_4787[40] ;
    input \prev_key1_new_127__N_4787[41] ;
    input \prev_key1_new_127__N_4787[42] ;
    input \prev_key1_new_127__N_4787[43] ;
    input \prev_key1_new_127__N_4787[44] ;
    input \prev_key1_new_127__N_4787[45] ;
    input \prev_key1_new_127__N_4787[46] ;
    input \prev_key1_new_127__N_4787[47] ;
    input \prev_key1_new_127__N_4787[48] ;
    input \prev_key1_new_127__N_4787[49] ;
    input \prev_key1_new_127__N_4787[50] ;
    input \prev_key1_new_127__N_4787[51] ;
    input \prev_key1_new_127__N_4787[52] ;
    input \prev_key1_new_127__N_4787[53] ;
    input \prev_key1_new_127__N_4787[54] ;
    input \prev_key1_new_127__N_4787[55] ;
    input \prev_key1_new_127__N_4787[56] ;
    input \prev_key1_new_127__N_4787[57] ;
    input \prev_key1_new_127__N_4787[58] ;
    input \prev_key1_new_127__N_4787[59] ;
    input \prev_key1_new_127__N_4787[60] ;
    input \prev_key1_new_127__N_4787[61] ;
    input \prev_key1_new_127__N_4787[62] ;
    input \prev_key1_new_127__N_4787[63] ;
    input n33431;
    input n33432;
    output n11_adj_123;
    input n33433;
    input n33434;
    input n33436;
    input n33441;
    input n33446;
    input n33448;
    input n33449;
    input n33450;
    input n33451;
    input n33452;
    input n33453;
    input n33454;
    input n33455;
    input n33456;
    input n33457;
    input n33458;
    input n33459;
    input n33460;
    input n33461;
    output n11_adj_124;
    input n33462;
    input n33463;
    input n33336;
    input n33435;
    input n33437;
    input n33438;
    input n33439;
    input n33440;
    input n33442;
    input n33443;
    input n33444;
    input n33445;
    input n33447;
    input n33337;
    input n33338;
    input n33339;
    input n33340;
    input n33341;
    input n33342;
    input n33350;
    input n33355;
    input n33361;
    input n33367;
    input n33374;
    input n33377;
    input n33379;
    input n33380;
    input n33382;
    input n33384;
    input n33386;
    output n11_adj_125;
    input n33387;
    input n33389;
    input n33391;
    input n33393;
    input n33395;
    input n33398;
    input n33400;
    input n33402;
    input n33405;
    input n33406;
    input n33409;
    input n33411;
    input n33413;
    output n11_adj_126;
    input [31:0]n2531;
    input n8532;
    input n9616;
    input n9618;
    input n9620;
    input n9622;
    input n9624;
    input n9626;
    input n9628;
    input n9630;
    input n9632;
    input n9634;
    input n9636;
    input n9638;
    input n9640;
    input n9642;
    input n9644;
    input n9646;
    input n9648;
    input n9650;
    input n9652;
    input n9654;
    input n9656;
    input n9658;
    input n9660;
    input n9662;
    output n11_adj_127;
    input n9664;
    input n9666;
    input n9668;
    input n9670;
    input n9672;
    input n9674;
    input n9676;
    input \key_mem_ctrl_new_2__N_4928[0] ;
    input block_w3_we_N_1490;
    input block_w2_we_N_1489;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(41[33:36])
    wire [127:0]\key_mem[6] ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(75[17:24])
    wire [127:0]\key_mem[7] ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(75[17:24])
    
    wire n5_c, n8, n9, n30758;
    wire [127:0]prev_key1_reg;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(83[17:30])
    wire [127:0]key_mem_new_127__N_7264;
    wire [127:0]\key_mem[12] ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(75[17:24])
    wire [127:0]\key_mem[13] ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(75[17:24])
    
    wire n1, n2, n30763, n33613, n8777;
    wire [127:0]prev_key0_reg;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(79[17:30])
    
    wire clk_c_enable_54;
    wire [127:0]prev_key0_new_127__N_4659;
    wire [7:0]rcon_reg;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(101[15:23])
    
    wire rcon_we;
    wire [7:0]rcon_new;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(102[15:23])
    
    wire n33614, n8775;
    wire [127:0]\key_mem[10] ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(75[17:24])
    wire [127:0]\key_mem[11] ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(75[17:24])
    
    wire n9_adj_8229;
    wire [127:0]\key_mem[8] ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(75[17:24])
    wire [127:0]\key_mem[9] ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(75[17:24])
    
    wire n8_adj_8230, n4, n33647;
    wire [7:0]\rcon_logic.tmp_rcon ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(314[19:27])
    
    wire n33716, n5_adj_8231;
    wire [127:0]\key_mem[4] ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(75[17:24])
    wire [127:0]\key_mem[5] ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(75[17:24])
    
    wire n4_adj_8232;
    wire [127:0]\key_mem[2] ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(75[17:24])
    wire [127:0]\key_mem[3] ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(75[17:24])
    
    wire n2_adj_8233;
    wire [127:0]\key_mem[0] ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(75[17:24])
    wire [127:0]\key_mem[1] ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(75[17:24])
    
    wire n1_adj_8234, n33717, n21, n21_adj_8235, n21_adj_8236, n21_adj_8237, 
        n21_adj_8238, n21_adj_8239, n21_adj_8240, n21_adj_8241, n21_adj_8242, 
        n21_adj_8243, n21_adj_8244, n21_adj_8245, n21_adj_8246, n21_adj_8247, 
        n21_adj_8248, n21_adj_8249, n21_adj_8250, n21_adj_8251, n21_adj_8252, 
        n21_adj_8253, n21_adj_8254, n21_adj_8255, n21_adj_8256, n21_adj_8257, 
        n21_adj_8258, n21_adj_8259, n21_adj_8260, n21_adj_8261, n21_adj_8262, 
        n21_adj_8263, n21_adj_8264, n22, n22_adj_8265, n22_adj_8266, 
        n22_adj_8267, n22_adj_8268, n22_adj_8269, n22_adj_8270, n22_adj_8271, 
        n22_adj_8272, n22_adj_8273, n22_adj_8274, n22_adj_8275, n22_adj_8276, 
        n22_adj_8277, n22_adj_8278, n22_adj_8279, n22_adj_8280, n22_adj_8281, 
        n22_adj_8282, n22_adj_8283, n22_adj_8284, n22_adj_8285, n22_adj_8286, 
        n22_adj_8287, n22_adj_8288, n22_adj_8289, n22_adj_8290, n22_adj_8291, 
        n33943, n33944, n28850, clk_c_enable_2335, n22_adj_8292, n22_adj_8293, 
        n22_adj_8294, n22_adj_8295;
    wire [127:0]n8680;
    
    wire clk_c_enable_2385, n9_adj_8308, n33718, n33859, n33547, n8_adj_8315, 
        n33615, n5_adj_8316, n4_adj_8317, n33719, n33616, n33738;
    wire [31:0]keymem_sboxw;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(107[18:30])
    
    wire n15897, n35839, n72, n2_adj_8318, n33747, n15304, n33720, 
        n1_adj_8319, n9_adj_8321, n8_adj_8322, n5_adj_8323, n4_adj_8324, 
        n2_adj_8325, n1_adj_8326, n2_adj_8328, n9_adj_8329, n8_adj_8330, 
        n33667, n15314, n33666, n35834, n8487, n1_adj_8331, n33664, 
        n15427, n33665, n8929, n33662, n15487, n33663, n4_adj_8332, 
        n33660, n15547, n33661, n4_adj_8333, n33658, n15607, n33659, 
        n4_adj_8335, n33656, n15667, n33657, n4_adj_8336, n33654, 
        n15727, n33655, n4_adj_8337, n33652, n15787, n33653, n9_adj_8338, 
        n4_adj_8339, n8_adj_8340, n33617, n33650, n15847, n33651, 
        n5_adj_8341, n4_adj_8342, n4_adj_8343, n2_adj_8344, n1_adj_8345, 
        n33648, n15907, n33649, n9_adj_8348, n4_adj_8349, n8_adj_8350, 
        n5_adj_8351, n9_adj_8352, n33646, n15967, n8_adj_8353, n4_adj_8354, 
        n5_adj_8355, n5_adj_8356, n4_adj_8357, n2_adj_8358, n4_adj_8359, 
        n33644, n16027, n33721, n33548, n33618, n33645, n1_adj_8360, 
        n4_adj_8361, n33722, n2_adj_8362, n33642, n16087, n9_adj_8364, 
        n33643, n2_adj_8365, n8_adj_8366, n4_adj_8367, n5_adj_8368, 
        n1_adj_8369, n4_adj_8370, n33640, n16147, n33641, n2_adj_8371, 
        n1_adj_8372, n4_adj_8373, n33638, n16207, n33639, n9_adj_8375, 
        n8_adj_8376, n4_adj_8377, n5_adj_8378, n33636, n16267, n4_adj_8379, 
        n33637, n2_adj_8380, n4_adj_8381, n1_adj_8382, n33634, n16327, 
        n1_adj_8383, n33723, n33619, n33635, n9_adj_8385, n4_adj_8386, 
        n8_adj_8387, n5_adj_8388, n33632, n16387, n33724, n33633, 
        n4_adj_8389, n4_adj_8390, n2_adj_8392, n1_adj_8393, n33630, 
        n16447, n33631, n4_adj_8395, n9_adj_8396, n8_adj_8397, n33628, 
        n16507, n33620, n33629, n5_adj_8398, clk_c_enable_104, n4_adj_8399, 
        n4_adj_8400, n2_adj_8401, n33626, n16567, n1_adj_8402, n33627, 
        n4_adj_8403, n9_adj_8404, n33624, n16627, n9_adj_8407, n33625, 
        n8_adj_8408, n8_adj_8409, n4_adj_8410, n5_adj_8411, n4_adj_8412, 
        n33622, n16687, n5_adj_8413, n2_adj_8414, n33623, n1_adj_8415, 
        n4_adj_8416, n4_adj_8417, n16747, n33621, n9_adj_8419, n8_adj_8420, 
        n4_adj_8421, n2_adj_8422, n5_adj_8423, n33572, n16807, n4_adj_8424, 
        n33573, n1_adj_8425, n2_adj_8426, n1_adj_8427, n4_adj_8428, 
        n33570, n16867, n33571;
    wire [31:0]\round_key_gen.trw ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(191[39:42])
    
    wire n4_adj_8430, n9_adj_8432, n8_adj_8433, n5_adj_8434, n4_adj_8435, 
        n33569, n16927, n33568, n9_adj_8436, n2_adj_8437, n4_adj_8438, 
        n1_adj_8439, n8_adj_8440, n33566, n16987, n33567, n9_adj_8442, 
        n8_adj_8443, n4_adj_8444, n5_adj_8445, n5_adj_8446, n4_adj_8447, 
        n4_adj_8448, n33564, n17047, n33565, n4_adj_8449, n2_adj_8450, 
        n33563, n17107, n33562, n4_adj_8451, n1_adj_8452, n33560, 
        n17167, n33561, n9_adj_8454, n4_adj_8455, n33559, n17227, 
        n33558, n8_adj_8456, n15124, n4_adj_8457, n5_adj_8458, n4_adj_8459, 
        n8711;
    wire [127:0]key_mem_new;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(76[17:28])
    
    wire n33557, n8713, n33746, n33556, n8715, n33745, n33555, 
        n8717, n2_adj_8460, n33744, n33554, n8719, n33743, n33553, 
        n8721, n33742, n33552, n9_adj_8461, n33739, n15837, n33725, 
        n1_adj_8462, n8723, n33741, n33551, n8725, n33740, n33550, 
        n8727, n33549, n8729, n8731, n9_adj_8464, n33737, n8733, 
        n8_adj_8465, n33736, n33546, n8735, n5_adj_8466, n8_adj_8467, 
        n33735, n33545, n4_adj_8468, n8737, n33734, n33544, n8739, 
        n2_adj_8469, n33733, n33543, n1_adj_8470, n33726, n5_adj_8471, 
        n8741, n33732, n33542, n4_adj_8472, n2_adj_8473, n8743, 
        n33731, n33541, n8745, n33730, n33540, n9_adj_8475, n1_adj_8476, 
        n8747, n8_adj_8477, n33729, n33539, n8749, n33728, n33538, 
        n5_adj_8478, n4_adj_8479, n8751, n33727, n33537, n2_adj_8480, 
        n8753, n33536, n1_adj_8481, n8755, n33535, n8757;
    wire [127:0]prev_key1_new_127__N_7520;
    
    wire n33534, n8759, n33517, n9_adj_8483, n8761, n8_adj_8484, 
        n8763, n33515, n5_adj_8485, n4_adj_8486, n8765, n33514, 
        n8767, n2_adj_8487, n33513, n1_adj_8488, n8769, n33512, 
        n8771, n8773, n9_adj_8491, n8_adj_8492, n5_adj_8493, n4_adj_8494, 
        n8779, n2_adj_8495, n1_adj_8496, n8781, n8783, n8785, n8787, 
        n8789, n9_adj_8498, n8791, n8_adj_8499, n8793, n5_adj_8500, 
        n4_adj_8501, n9_adj_8502, n8795, n8797, n2_adj_8503, n8799, 
        n1_adj_8504, n8801, n8803, n8805, n9_adj_8506, n8807, n8809, 
        n8_adj_8507, n8811, n8_adj_8508, n5_adj_8509, n4_adj_8510, 
        n8813, n2_adj_8511, n8815, n8817, n1_adj_8512, n8819, n8821, 
        n8823, n8825, n9_adj_8514, n33532, n8_adj_8515, n8827, n8829, 
        n8831, n5_adj_8516, n4_adj_8517, n8833, n2_adj_8518, n8835, 
        n33527, n8837, n33526, n1_adj_8519, n9_adj_8521, n8_adj_8522, 
        n5_adj_8523, n4_adj_8524, n2_adj_8525, n1_adj_8526, n9_adj_8528, 
        n8_adj_8529, n5_adj_8530, n4_adj_8531, n2_adj_8532, n1_adj_8533, 
        n5_adj_8535, n4_adj_8536, n9_adj_8537, n8_adj_8538, n5_adj_8539, 
        n4_adj_8540, n2_adj_8541, n15777, n2_adj_8542, n1_adj_8543, 
        n1_adj_8545, n9_adj_8546, n8_adj_8547, n9_adj_8549, n8_adj_8550, 
        n5_adj_8551, n4_adj_8552, n2_adj_8553, n1_adj_8554, n5_adj_8555, 
        n9_adj_8557, n8_adj_8558, n5_adj_8559, n4_adj_8560, n4_adj_8561, 
        n2_adj_8562, n1_adj_8563, clk_c_enable_436;
    wire [127:0]key_mem_0__127__N_6752;
    wire [127:0]prev_key1_new_127__N_4787;
    
    wire n2_adj_8565, n1_adj_8566, n9_adj_8567, n8_adj_8568, n10;
    wire [31:0]muxed_sboxw;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(109[18:29])
    
    wire n9_adj_8571, n8_adj_8572, n5_adj_8573, n4_adj_8574, n15717, 
        n2_adj_8575, n1_adj_8576, n5_adj_8577, n9_adj_8579, n8_adj_8580, 
        n4_adj_8581, n5_adj_8582, n4_adj_8583, n2_adj_8584, n1_adj_8585, 
        n10_adj_8587, n2_adj_8588, n1_adj_8589, n10_adj_8590, n9_adj_8591, 
        n8_adj_8592, n5_adj_8593, n4_adj_8594, n2_adj_8595, n1_adj_8597, 
        n10_adj_8598, n9_adj_8599, n8_adj_8601, n10_adj_8602, n5_adj_8603, 
        n4_adj_8604, n15657, n9_adj_8605, n8_adj_8606, n10_adj_8607, 
        n10_adj_8608, n5_adj_8609, n4_adj_8610, n2_adj_8611, n2_adj_8612, 
        n1_adj_8613, n10_adj_8614, n10_adj_8615, n1_adj_8616, n10_adj_8617, 
        n9_adj_8619, n10_adj_8620, n8_adj_8621, n10_adj_8622, n5_adj_8623, 
        n4_adj_8624, n10_adj_8625, n10_adj_8627, n2_adj_8628, n1_adj_8629, 
        n9_adj_8631, n8_adj_8632, n10_adj_8633, n5_adj_8634, n4_adj_8635, 
        n9_adj_8636, n10_adj_8637, n2_adj_8638, n10_adj_8639, n10_adj_8640, 
        n8_adj_8641, n10_adj_8642, n1_adj_8643, n10_adj_8644, n10_adj_8645, 
        n5_adj_8646, n10_adj_8648, n4_adj_8649, n10_adj_8650, n10_adj_8651, 
        n9_adj_8652, n8_adj_8653, n5_adj_8654, n4_adj_8655, n2_adj_8656, 
        n1_adj_8657, n8478, n2958;
    wire [3:0]n6361;
    
    wire n33951, key_mem_ctrl_we, n7;
    wire [3:0]round_ctr_reg;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(87[15:28])
    
    wire n33912, n9_adj_8660, n9_adj_8661, n8_adj_8662, n8_adj_8663, 
        n5_adj_8664, n4_adj_8665, n5_adj_8666, n2_adj_8667, n4_adj_8668, 
        n1_adj_8669, n2_adj_8670, n9_adj_8672, n8_adj_8673, n1_adj_8674, 
        n2_adj_8675, n1_adj_8676, n15597, n5_adj_8677, n4_adj_8678, 
        n2_adj_8680, n9_adj_8681, n8_adj_8682, n1_adj_8683, n9_adj_8685, 
        n8_adj_8686, n5_adj_8687, n4_adj_8688, n15537, n15477, n2_adj_8689, 
        n15417, n1_adj_8690, n9_adj_8692, n8_adj_8693, n5_adj_8694, 
        n4_adj_8695, n2_adj_8696, n1_adj_8697, n9_adj_8699, n8_adj_8700, 
        n5_adj_8701, n4_adj_8702, n5_adj_8703, n4_adj_8705, n2_adj_8706, 
        n9_adj_8707, n1_adj_8708, n2_adj_8709, n30840, n8_adj_8710, 
        n5_adj_8711, n1_adj_8712, n4_adj_8713, n2_adj_8714, n1_adj_8715, 
        n9_adj_8717, n8_adj_8718, n5_adj_8719, n4_adj_8720, n9_adj_8722, 
        n8_adj_8723, n5_adj_8724, n4_adj_8725, n2_adj_8726, n2_adj_8727, 
        n1_adj_8728, n1_adj_8729, n9_adj_8732, n9_adj_8733, n8_adj_8734, 
        n8_adj_8735, n5_adj_8736, n5_adj_8737, n4_adj_8738, n4_adj_8739, 
        n2_adj_8740, n1_adj_8741, n2_adj_8742, n1_adj_8743, n9_adj_8746, 
        n8_adj_8747, n5_adj_8748, n9_adj_8749, n8_adj_8750, n4_adj_8751, 
        n5_adj_8752, n4_adj_8753, n2_adj_8754, n2_adj_8755, n1_adj_8756, 
        n1_adj_8757, n9_adj_8759, n8_adj_8760, n9_adj_8762, n5_adj_8763, 
        n4_adj_8764, n8_adj_8765, n2_adj_8766, n5_adj_8767, n1_adj_8768, 
        n4_adj_8769, n2_adj_8771, n1_adj_8772, n9_adj_8773, n8_adj_8774, 
        n5_adj_8776, n4_adj_8777, n2_adj_8778, n1_adj_8779, n9_adj_8780, 
        n8_adj_8781, n5_adj_8782, n4_adj_8783, n2_adj_8785, n1_adj_8786, 
        n9_adj_8787, n8_adj_8788, n5_adj_8789, n4_adj_8791, n2_adj_8792, 
        n1_adj_8793, n9_adj_8794, n8_adj_8795, n9_adj_8797, n5_adj_8798, 
        n8_adj_8799, n5_adj_8800, n4_adj_8801, n4_adj_8802, n2_adj_8803, 
        n2_adj_8804, n1_adj_8805, n1_adj_8806, n9_adj_8808, n8_adj_8809, 
        n5_adj_8811, n4_adj_8812, n2_adj_8813, n9_adj_8814, n1_adj_8815, 
        n8_adj_8816, n5_adj_8818, n9_adj_8819, n8_adj_8820, n4_adj_8821, 
        n2_adj_8822, n5_adj_8823, n1_adj_8824, n4_adj_8825, n2_adj_8826, 
        n1_adj_8827, n9_adj_8830, n8_adj_8831, n9_adj_8832, n8_adj_8833, 
        n5_adj_8834, n5_adj_8835, n4_adj_8836, n4_adj_8837, n2_adj_8838, 
        n2_adj_8839, n1_adj_8840, n1_adj_8841, n9_adj_8843, n8_adj_8845, 
        n9_adj_8846, n5_adj_8847, n4_adj_8848, n8_adj_8849, n2_adj_8850, 
        n1_adj_8851, n5_adj_8852, n4_adj_8853, n9_adj_8855, n2_adj_8856, 
        n8_adj_8857, n1_adj_8858, n5_adj_8859, n4_adj_8860, n2_adj_8861, 
        n1_adj_8863, n9_adj_8864, n8_adj_8866, n9_adj_8867, n8_adj_8868, 
        n5_adj_8869, n5_adj_8870, n4_adj_8871, n4_adj_8872, n2_adj_8873, 
        n1_adj_8874, n2_adj_8875, n1_adj_8876, n9_adj_8878, n8_adj_8879, 
        n5_adj_8881, n4_adj_8882, n9_adj_8883, n2_adj_8884, n1_adj_8885, 
        n8_adj_8886, n5_adj_8888, n4_adj_8889, n9_adj_8890, n2_adj_8891, 
        n8_adj_8892, n1_adj_8893, n5_adj_8894, n4_adj_8895, n33528, 
        n2_adj_8897, n30151, n30152, n9_adj_8898, n1_adj_8899, n30158, 
        n30159, n8_adj_8900, n30165, n30166, n5_adj_8902, n4_adj_8903, 
        n9_adj_8904, n2_adj_8905, n8_adj_8906, n1_adj_8907, n5_adj_8908, 
        n4_adj_8909, n33510, n30172, n30173, n2_adj_8910, n1_adj_8911, 
        n30179, n30180, n33529, n9_adj_8914, n9_adj_8915, n8_adj_8916, 
        n8_adj_8917, n5_adj_8918, n4_adj_8919, n5_adj_8920, n4_adj_8922, 
        n33530, n9_adj_8923, n30186, n30187, n8_adj_8924, n2_adj_8925, 
        n1_adj_8926, n5_adj_8927, n4_adj_8928, n30193, n30194, n30200, 
        n30201, n2_adj_8930, n1_adj_8931, n9_adj_8932, n8_adj_8933, 
        n5_adj_8934, n33531, n4_adj_8936, n30207, n30208, n2_adj_8937, 
        n1_adj_8938, n30214, n30215, n9_adj_8940, n9_adj_8941, n30221, 
        n30222, n30228, n30229, n8_adj_8942, n30235, n30236, n30242, 
        n30243, n5_adj_8943, n30249, n30250, n30256, n30257, n4_adj_8944, 
        n2_adj_8945, n1_adj_8946, n8_adj_8947, n30263, n30264, n30270, 
        n30271, n30277, n30278, n33533, n9_adj_8949, n8_adj_8950, 
        n30284, n30285, n5_adj_8951, n5_adj_8952, n4_adj_8953, n4_adj_8954, 
        n30291, n30292, n30298, n30299, n30305, n30306, n30312, 
        n30313, n30319, n30320, n30326, n30327, n2_adj_8955, n4_adj_8956, 
        n5_adj_8957, n30841, n30333, n30334, n1_adj_8958, n33511, 
        n2_adj_8959, n30340, n30341, n1_adj_8960, n30347, n30348, 
        n9_adj_8962, n30354, n30355, n30361, n30362, n30368, n30369, 
        n30375, n30376, n8_adj_8963, n30382, n30383, n5_adj_8964, 
        n30389, n30390, n30396, n30397, n4_adj_8965, n30403, n30404, 
        n2_adj_8966, n30410, n30411, n30417, n30418, n1_adj_8967, 
        n30424, n30425, n30431, n30432, n30438, n30439, n30445, 
        n30446, n30452, n30453, n30459, n30460, n30466, n30467, 
        n9_adj_8970, n30473, n30474, n30480, n30481, n8_adj_8971, 
        n5_adj_8972, n30487, n30488, n30494, n30495, n30501, n30502, 
        n4_adj_8973, n2_adj_8974, n1_adj_8975, n9_adj_8976, n8_adj_8977, 
        n9_adj_8979, n4_adj_8980, n16742, n8_adj_8981, n5_adj_8982, 
        n4_adj_8983, n4_adj_8984, n16682, n2_adj_8985, n5_adj_8986, 
        n1_adj_8987, n4_adj_8988, n16622, n4_adj_8990, n16562, n4_adj_8991, 
        n9_adj_8992, n4_adj_8993, n16502, n8_adj_8994, n4_adj_8995, 
        n16442, n5_adj_8996, n4_adj_8997, n2_adj_8998, n1_adj_8999, 
        n4_adj_9000, n16382, n4_adj_9001, n16322, n2_adj_9002, n17097, 
        n4_adj_9003, n16262, n1_adj_9005, n9_adj_9006, n4_adj_9007, 
        n16202, n8_adj_9008, n5_adj_9009, n4_adj_9010, n4_adj_9011, 
        n16142, n2_adj_9012, n4_adj_9013, n16082, n1_adj_9014, n17037, 
        n4_adj_9015, n16022, n9_adj_9017, n8_adj_9018, n4_adj_9019, 
        n15962, n30508, n30509, n30515, n30516, n4_adj_9021, n15902, 
        n5_adj_9022, n4_adj_9023, n4_adj_9024, n15842, n2_adj_9025, 
        n30522, n30523, n30529, n30530, n30536, n30537, n30543, 
        n30544, n30550, n30551, n30557, n30558, n30564, n30565, 
        n30571, n30572, n30578, n30579, n30585, n30586, n30592, 
        n30593, n1_adj_9026, n4_adj_9027, n15782, n30599, n30600, 
        n30606, n30607, n30613, n30614, n30620, n30621, n4_adj_9029, 
        n15722, n30627, n30628, n9_adj_9030, n30634, n30635, n8_adj_9031, 
        n30641, n30642, n30648, n30649, n30655, n30656, n30662, 
        n30663, n30669, n30670, n30676, n30677, n30683, n30684, 
        n30690, n30691, n30697, n30698, n30704, n30705, n30711, 
        n30712, n4_adj_9032, n15662, n30718, n30719, n30725, n30726, 
        n30732, n30733, n5_adj_9033, n30739, n30740, n30746, n30747, 
        n30753, n30754, n30760, n30761, n30767, n30768, n30774, 
        n30775, n30781, n30782, n30788, n30789, n30795, n30796, 
        n30802, n30803, n30809, n30810, n4_adj_9034, n15602, n30816, 
        n30817, n30823, n30824, n30830, n30831, n4_adj_9035, n30837, 
        n30838, n9_adj_9036, n30844, n30845, n8_adj_9037, n30851, 
        n30852, n30858, n30859, n30865, n30866, n2_adj_9038, n30872, 
        n30873, n30879, n30880, n1_adj_9039, n30886, n30887, n30893, 
        n30894, n30900, n30901, n30907, n30908, n30914, n30915, 
        n30921, n30922, n4_adj_9040, n15542, n31024, n31025, n31031, 
        n31032, n31038, n31039, n31045, n31046, n31052, n31053, 
        n31059, n31060, n31066, n31067, n31073, n31074, n31080, 
        n31081, n31087, n31088, n31094, n31095, n31101, n31102, 
        n31108, n31109, n31115, n31116, n31122, n31123, n31129, 
        n31130, n31136, n31137, n30147, n30148, n4_adj_9042, n15482, 
        n30149, n9_adj_9043, n5_adj_9044, n30154, n30155, n30156, 
        n30161, n30162, n30163, n4_adj_9045, n30168, n30169, n30170, 
        n4_adj_9046, n15422, n30175, n30176, n30177, n30182, n30183, 
        n30184, n30189, n30190, n30191, n30196, n30197, n30198, 
        n30203, n30204, n30205, n30210, n30211, n30212, n30217, 
        n30218, n30219, n30224, n30225, n30226, n30231, n30232, 
        n30233, n30238, n30239, n8_adj_9047, n30240, n30245, n30246, 
        n4_adj_9048, n15309, n30247, n5_adj_9049, n4_adj_9050, n30252, 
        n30253, n4_adj_9051, n17222, n2_adj_9052, n30254, n1_adj_9053, 
        n30259, n30260, n30261, n30266, n30267, n30268, n30273, 
        n30274, n30275, n30280, n30281, n30282, n30287, n30288, 
        n4_adj_9054, n17162, n4_adj_9055, n17102, n9_adj_9057, n8_adj_9058, 
        n4_adj_9059, n17042, n5_adj_9060, n4_adj_9061, n16982, n30289, 
        n30294, n30295, n30296, n30301, n30302, n30303, n30308, 
        n30309, n30310, n4_adj_9062, n30315, n30316, n30317, n30322, 
        n30323, n2_adj_9063, n4_adj_9064, n16922, n1_adj_9065, n4_adj_9067, 
        n16862, n9_adj_9068, n30324, n30329, n30330, n30331, n30336, 
        n30337, n30338, n8_adj_9069, n30343, n30344, n30345, n15311, 
        n30350, n30351, n30352, n30357, n30358, n5_adj_9070, n30359, 
        n4_adj_9071, n30364, n30365, n2_adj_9072, n30366, n1_adj_9073, 
        n30371, n30372, n30373, n30378, n30379, n30380, n30385, 
        n30386, n30387, n30392, n30393, n16977, n9_adj_9075, n8_adj_9076, 
        n5_adj_9077, n2_adj_9078, n4_adj_9079, n1_adj_9080, n2_adj_9081, 
        n1_adj_9082, n4_adj_9084, n16802, n9_adj_9085, n8_adj_9086, 
        n5_adj_9087, n4_adj_9088, n2_adj_9089, n30394, n1_adj_9091, 
        n9_adj_9092, n8_adj_9093, n9_adj_9095, n8_adj_9096, n5_adj_9097, 
        n4_adj_9098, n2_adj_9099, n1_adj_9100, n9_adj_9102, n8_adj_9103, 
        n5_adj_9104, n4_adj_9105, n2_adj_9106, n1_adj_9107, n9_adj_9109, 
        n8_adj_9110, n5_adj_9111, n4_adj_9112, n2_adj_9113, n1_adj_9114, 
        n5_adj_9115, n4_adj_9116, n9_adj_9118, n2_adj_9119, n1_adj_9120, 
        n8_adj_9121, n33911, n5_adj_9123, n9_adj_9124, n4_adj_9125, 
        n2_adj_9126, n8_adj_9127, n1_adj_9128, n5_adj_9129, n16917, 
        n9_adj_9131, n8_adj_9132, n5_adj_9133, n4_adj_9134, n2_adj_9135, 
        n1_adj_9136, n4_adj_9137, n9_adj_9139, n8_adj_9140, n5_adj_9141, 
        n4_adj_9142, n2_adj_9143, n1_adj_9144, n2_adj_9145, n9_adj_9147, 
        n8_adj_9148, n5_adj_9149, n4_adj_9150, n1_adj_9151, n2_adj_9152, 
        n1_adj_9153, n9_adj_9156, n8_adj_9157, n5_adj_9158, n4_adj_9159, 
        n2_adj_9160, n1_adj_9161, n33516, n9_adj_9163, n9_adj_9164, 
        n8_adj_9165, n30399, n30400, n30401, n5_adj_9166, n4_adj_9167, 
        n2_adj_9168, n1_adj_9169, n9_adj_9171, n30406, n30407, n30408, 
        n8_adj_9172, n30413, n30414, n5_adj_9173, n30415, n4_adj_9174, 
        n30420, n30421, n2_adj_9175, n30422, n1_adj_9176, n30427, 
        n30428, n16797, n30429, n30434, n30435, n30436, n30441, 
        n30442, n9_adj_9178, n8_adj_9179, n5_adj_9180, n4_adj_9181, 
        n2_adj_9182, n1_adj_9183, n9_adj_9185, n8_adj_9186, n5_adj_9187, 
        n4_adj_9188, n2_adj_9189, n1_adj_9190, n9_adj_9192, n8_adj_9193, 
        n5_adj_9194, clk_c_enable_132, n30443, n4_adj_9195, n30448, 
        n30449, n2_adj_9196, n30450, n1_adj_9197, n30455, n30456, 
        n30457, n30462, n30463, n30464, n30469, n30470, n9_adj_9199, 
        n8_adj_9200, n30471, n5_adj_9201, n4_adj_9202, n30476, n30477, 
        n30478, n30483, n30484, n2_adj_9203, n30485, n1_adj_9204, 
        n30490, n30491, n8_adj_9205, n30492, n30497, n30498, n9_adj_9207, 
        n30499, n8_adj_9208, n30504, n30505, n5_adj_9209, n4_adj_9210, 
        n30506, n2_adj_9211, n30511, n30512, n1_adj_9212, n30513, 
        n2_adj_9213, n30518, n30519, n1_adj_9214, n30520, n30525, 
        n30526, n30527, n30532, n30533, n5_adj_9215, n30534, n30539, 
        n30540, n30541, n30546, n30547, n30548, n30553, n30554, 
        n4_adj_9216, n30555, n30560, n30561, n30562, n30567, n30568, 
        n4_adj_9217, n30569, n30574, n30575, n30576, n2_adj_9218, 
        n1_adj_9219, n30581, n30582, n30583, n30588, n30589, n30590, 
        n30595, n30596;
    wire [127:0]key_mem_0__127__N_5216;
    
    wire n2_adj_9220, n1_adj_9221, n9_adj_9223, n8_adj_9224, n5_adj_9225, 
        n4_adj_9226, n2_adj_9227, n1_adj_9228, n9_adj_9230, n8_adj_9231, 
        n5_adj_9232, n4_adj_9233, n2_adj_9234, n1_adj_9235, n9_adj_9237, 
        n8_adj_9238, n5_adj_9239, n4_adj_9240, n2_adj_9241, n1_adj_9242, 
        n9_adj_9244, n8_adj_9245, n5_adj_9246, n4_adj_9247, n2_adj_9248, 
        n1_adj_9249, n9_adj_9251, n8_adj_9252, n33938;
    wire [127:0]key_mem_0__127__N_5344;
    
    wire clk_c_enable_486, clk_c_enable_536;
    wire [127:0]key_mem_0__127__N_6624;
    
    wire clk_c_enable_586, clk_c_enable_636, clk_c_enable_686;
    wire [127:0]key_mem_0__127__N_6496;
    
    wire clk_c_enable_736, clk_c_enable_786;
    wire [127:0]key_mem_0__127__N_6368;
    
    wire clk_c_enable_836, clk_c_enable_886, clk_c_enable_936;
    wire [127:0]key_mem_0__127__N_6240;
    
    wire clk_c_enable_986, clk_c_enable_1036;
    wire [127:0]key_mem_0__127__N_6112;
    
    wire clk_c_enable_1086, clk_c_enable_1136, clk_c_enable_1186;
    wire [127:0]key_mem_0__127__N_5984;
    
    wire clk_c_enable_1236, clk_c_enable_1286;
    wire [127:0]key_mem_0__127__N_5856;
    
    wire clk_c_enable_1336, clk_c_enable_1386, clk_c_enable_1436;
    wire [127:0]key_mem_0__127__N_5728;
    
    wire clk_c_enable_1486, clk_c_enable_1536, clk_c_enable_1586;
    wire [127:0]key_mem_0__127__N_5600;
    
    wire clk_c_enable_1636, clk_c_enable_1686;
    wire [127:0]key_mem_0__127__N_5472;
    
    wire clk_c_enable_1736, clk_c_enable_1786, clk_c_enable_1836, clk_c_enable_1886, 
        clk_c_enable_1936, clk_c_enable_1986, clk_c_enable_2036, clk_c_enable_2086;
    wire [127:0]key_mem_0__127__N_5088;
    
    wire clk_c_enable_2136, clk_c_enable_2186;
    wire [127:0]key_mem_0__127__N_4960;
    
    wire clk_c_enable_2236, clk_c_enable_2286, clk_c_enable_2413, n30597, 
        n30602, n30603, n30604, n30609, n30610, n30611, n30616, 
        n30617, n30618, n9_adj_9254, n8_adj_9255, n30623, n30624, 
        n30625, n30630, n30631, n30632, n10_adj_9256, n30637, n30638, 
        n5_adj_9257, n30639, n30644, n30645, n30646, n10_adj_9258, 
        n4_adj_9259, n30651, n30652, n30653, n30658, n30659, n10_adj_9260, 
        n30660, n10_adj_9261, n30665, n30666, n30667, n2_adj_9262, 
        n30672, n30673, n1_adj_9263, n30674, n30679, n30680, n30842, 
        n30681, n33591, n30686, n30687, n30688, n30847, n30693, 
        n30694, n33592, n30695, n30700, n30701, n30848, n30702, 
        n30707, n30708, n30709, n10_adj_9264, n30849, n30714, n30715, 
        n30716, n30721, n30722, n30723, n33593, n30728, n30729, 
        n30730, n30854, n30735, n30736, n30737, n30855, n30742, 
        n30743, n30744, n33594, n30749, n30750, n30751, n30756, 
        n30757, n30764, n30856, n30765, n30770, n30771, n30772, 
        n33595, n9_adj_9266, n30777, n30778, n30779, n8_adj_9267, 
        n10_adj_9268, n30784, n30785, n30786, n30861, n33596, n30791, 
        n30792, n30793, n30862, n30798, n30799, n30800, n30863, 
        n33597, n30805, n30806, n5_adj_9269, n30807, n30812, n30813, 
        n10_adj_9270, n30814, n4_adj_9271, n10_adj_9272, n30819, n30820, 
        n30821, n30826, n30827, n30828, n30868, n30833, n30834, 
        n33598, n30835, n30869, n2_adj_9273, n30870, n33599, n33916, 
        n1_adj_9274, n30875, n30876, n30877, n33600, n30882, n30883, 
        n30884, n16017, n30889, n30890, n30891, n30896, n30897, 
        n30898, n33601, n30903, n30904, n30905, n30910, n30911, 
        n30912, n30917, n30918, n30919, n31020, n31021, n33602, 
        n31022, n31027, n31028, n31029, n33603, n33945, n31034, 
        n31035, n31036, n31041, n31042, n31043, n31048, n31049, 
        n31050, n31055, n31056, n31057, n33604, n31062, n31063, 
        n31064, n31069, n31070, n31071, n33605, n31076, n31077, 
        n31078, n31083, n31084, n31085, n31090, n31091, n31092, 
        n9_adj_9276, n31097, n31098, n31099, n8_adj_9277, n31104, 
        n31105, n31106, n31111, n31112, n31113, n33606, n31118, 
        n31119, n31120, n5_adj_9278, n4_adj_9279, n31125, n31126, 
        n31127, n33607, n31132, n31133, n31134, n2_adj_9280, n33608, 
        n1_adj_9281, n33609, n33610, n9_adj_9283, n8_adj_9284, n5_adj_9285, 
        n33611, n15957, n4_adj_9286, n2_adj_9287, n33612, n1_adj_9288, 
        round_ctr_we;
    wire [3:0]n3;
    
    wire n15086, n1_adj_9290, n33937, n16803, n16857, n16863, n16923, 
        n16983, n17043, n17103, n17157, n17163, n17217, n17223, 
        n15310, n15423, n15483, n15543, n15603, n15663, n15723, 
        n15783, n15843, n15903, n15963, n16023, n16077, n16083, 
        n16137, n16143, n16197, n16203, n16257, n16263, n16317, 
        n16323, n16377, n16383, n16437, n16443, n16497, n16503, 
        n16557, n16563, n16617, n16623, n16677, n16683, n16737, 
        n16743, n28834, n29504, n21_adj_9291, n2952;
    
    LUT4 round_3__I_0_Mux_104_i5_3_lut (.A(\key_mem[6] [104]), .B(\key_mem[7] [104]), 
         .C(n33952), .Z(n5_c)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_104_i5_3_lut.init = 16'hcaca;
    PFUMX i25599 (.BLUT(n8), .ALUT(n9), .C0(\muxed_round_nr[1] ), .Z(n30758));
    LUT4 mux_51_i99_3_lut_4_lut (.A(prev_key1_reg[98]), .B(\round_key_gen.trw[2] ), 
         .C(n33860), .D(\key_reg[0] [2]), .Z(key_mem_new_127__N_7264[98])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam mux_51_i99_3_lut_4_lut.init = 16'h6f60;
    LUT4 round_3__I_0_Mux_99_i11_3_lut (.A(\key_mem[12] [99]), .B(\key_mem[13] [99]), 
         .C(n33952), .Z(n11)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_99_i11_3_lut.init = 16'hcaca;
    PFUMX i25604 (.BLUT(n1), .ALUT(n2), .C0(\muxed_round_nr[1] ), .Z(n30763));
    LUT4 i3292_3_lut_4_lut (.A(prev_key1_reg[97]), .B(\round_key_gen.trw[1] ), 
         .C(n35835), .D(n33613), .Z(n8777)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam i3292_3_lut_4_lut.init = 16'hf606;
    FD1P3IX prev_key0_reg__i0 (.D(prev_key0_new_127__N_4659[0]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i0.GSR = "DISABLED";
    LUT4 mux_51_i98_3_lut_4_lut (.A(prev_key1_reg[97]), .B(\round_key_gen.trw[1] ), 
         .C(n33860), .D(\key_reg[0] [1]), .Z(key_mem_new_127__N_7264[97])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam mux_51_i98_3_lut_4_lut.init = 16'h6f60;
    FD1P3AX rcon_reg_i0_i0 (.D(rcon_new[0]), .SP(rcon_we), .CK(clk_c), 
            .Q(rcon_reg[0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam rcon_reg_i0_i0.GSR = "ENABLED";
    LUT4 i3290_3_lut_4_lut (.A(prev_key1_reg[96]), .B(\round_key_gen.trw[0] ), 
         .C(n35835), .D(n33614), .Z(n8775)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam i3290_3_lut_4_lut.init = 16'hf606;
    LUT4 round_3__I_0_Mux_99_i9_3_lut (.A(\key_mem[10] [99]), .B(\key_mem[11] [99]), 
         .C(n33952), .Z(n9_adj_8229)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_99_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_99_i8_3_lut (.A(\key_mem[8] [99]), .B(\key_mem[9] [99]), 
         .C(n33952), .Z(n8_adj_8230)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_99_i8_3_lut.init = 16'hcaca;
    LUT4 i2_2_lut_rep_343 (.A(prev_key0_reg[74]), .B(n4), .Z(n33647)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i2_2_lut_rep_343.init = 16'h6666;
    LUT4 mux_51_i97_3_lut_4_lut (.A(prev_key1_reg[96]), .B(\round_key_gen.trw[0] ), 
         .C(n33860), .D(\key_reg[0] [0]), .Z(key_mem_new_127__N_7264[96])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam mux_51_i97_3_lut_4_lut.init = 16'h6f60;
    LUT4 i2_3_lut_rep_412 (.A(\new_sboxw[23] ), .B(\rcon_logic.tmp_rcon [0]), 
         .C(prev_key1_reg[127]), .Z(n33716)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(110[18:27])
    defparam i2_3_lut_rep_412.init = 16'h9696;
    LUT4 round_3__I_0_Mux_99_i5_3_lut (.A(\key_mem[6] [99]), .B(\key_mem[7] [99]), 
         .C(n33952), .Z(n5_adj_8231)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_99_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_99_i4_3_lut (.A(\key_mem[4] [99]), .B(\key_mem[5] [99]), 
         .C(n33952), .Z(n4_adj_8232)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_99_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_99_i2_3_lut (.A(\key_mem[2] [99]), .B(\key_mem[3] [99]), 
         .C(n33952), .Z(n2_adj_8233)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_99_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_99_i1_3_lut (.A(\key_mem[0] [99]), .B(\key_mem[1] [99]), 
         .C(n33952), .Z(n1_adj_8234)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_99_i1_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_rep_413 (.A(\new_sboxw[22] ), .B(prev_key1_reg[126]), 
         .C(\rcon_logic.tmp_rcon [7]), .Z(n33717)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(110[18:27])
    defparam i2_3_lut_rep_413.init = 16'h9696;
    LUT4 i1_4_lut (.A(\key_mem_ctrl.num_rounds[2] ), .B(\key_reg[3] [1]), 
         .C(n21), .D(n33860), .Z(prev_key0_new_127__N_4659[1])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(85[17:29])
    defparam i1_4_lut.init = 16'ha088;
    LUT4 i1_4_lut_adj_488 (.A(\key_mem_ctrl.num_rounds[2] ), .B(\key_reg[3] [2]), 
         .C(n21_adj_8235), .D(n33860), .Z(prev_key0_new_127__N_4659[2])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(85[17:29])
    defparam i1_4_lut_adj_488.init = 16'ha088;
    LUT4 i1_4_lut_adj_489 (.A(\key_mem_ctrl.num_rounds[2] ), .B(\key_reg[3] [3]), 
         .C(n21_adj_8236), .D(n33860), .Z(prev_key0_new_127__N_4659[3])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(85[17:29])
    defparam i1_4_lut_adj_489.init = 16'ha088;
    LUT4 i1_4_lut_adj_490 (.A(\key_mem_ctrl.num_rounds[2] ), .B(\key_reg[3] [4]), 
         .C(n21_adj_8237), .D(n33860), .Z(prev_key0_new_127__N_4659[4])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(85[17:29])
    defparam i1_4_lut_adj_490.init = 16'ha088;
    LUT4 i1_4_lut_adj_491 (.A(\key_mem_ctrl.num_rounds[2] ), .B(\key_reg[3] [5]), 
         .C(n21_adj_8238), .D(n33860), .Z(prev_key0_new_127__N_4659[5])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(85[17:29])
    defparam i1_4_lut_adj_491.init = 16'ha088;
    LUT4 i1_4_lut_adj_492 (.A(\key_mem_ctrl.num_rounds[2] ), .B(\key_reg[3] [6]), 
         .C(n21_adj_8239), .D(n33860), .Z(prev_key0_new_127__N_4659[6])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(85[17:29])
    defparam i1_4_lut_adj_492.init = 16'ha088;
    LUT4 i1_4_lut_adj_493 (.A(\key_mem_ctrl.num_rounds[2] ), .B(\key_reg[3] [7]), 
         .C(n21_adj_8240), .D(n33860), .Z(prev_key0_new_127__N_4659[7])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(85[17:29])
    defparam i1_4_lut_adj_493.init = 16'ha088;
    LUT4 i1_4_lut_adj_494 (.A(\key_mem_ctrl.num_rounds[2] ), .B(\key_reg[3] [8]), 
         .C(n21_adj_8241), .D(n33860), .Z(prev_key0_new_127__N_4659[8])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(85[17:29])
    defparam i1_4_lut_adj_494.init = 16'ha088;
    LUT4 i1_4_lut_adj_495 (.A(\key_mem_ctrl.num_rounds[2] ), .B(\key_reg[3] [9]), 
         .C(n21_adj_8242), .D(n33860), .Z(prev_key0_new_127__N_4659[9])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(85[17:29])
    defparam i1_4_lut_adj_495.init = 16'ha088;
    LUT4 i1_4_lut_adj_496 (.A(\key_mem_ctrl.num_rounds[2] ), .B(\key_reg[3] [10]), 
         .C(n21_adj_8243), .D(n33860), .Z(prev_key0_new_127__N_4659[10])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(85[17:29])
    defparam i1_4_lut_adj_496.init = 16'ha088;
    LUT4 i1_4_lut_adj_497 (.A(\key_mem_ctrl.num_rounds[2] ), .B(\key_reg[3] [11]), 
         .C(n21_adj_8244), .D(n33860), .Z(prev_key0_new_127__N_4659[11])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(85[17:29])
    defparam i1_4_lut_adj_497.init = 16'ha088;
    LUT4 i1_4_lut_adj_498 (.A(\key_mem_ctrl.num_rounds[2] ), .B(\key_reg[3] [12]), 
         .C(n21_adj_8245), .D(n33860), .Z(prev_key0_new_127__N_4659[12])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(85[17:29])
    defparam i1_4_lut_adj_498.init = 16'ha088;
    LUT4 i1_4_lut_adj_499 (.A(\key_mem_ctrl.num_rounds[2] ), .B(\key_reg[3] [13]), 
         .C(n21_adj_8246), .D(n33860), .Z(prev_key0_new_127__N_4659[13])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(85[17:29])
    defparam i1_4_lut_adj_499.init = 16'ha088;
    LUT4 i1_4_lut_adj_500 (.A(\key_mem_ctrl.num_rounds[2] ), .B(\key_reg[3] [14]), 
         .C(n21_adj_8247), .D(n33860), .Z(prev_key0_new_127__N_4659[14])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(85[17:29])
    defparam i1_4_lut_adj_500.init = 16'ha088;
    LUT4 i1_4_lut_adj_501 (.A(\key_mem_ctrl.num_rounds[2] ), .B(\key_reg[3] [15]), 
         .C(n21_adj_8248), .D(n33860), .Z(prev_key0_new_127__N_4659[15])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(85[17:29])
    defparam i1_4_lut_adj_501.init = 16'ha088;
    LUT4 i1_4_lut_adj_502 (.A(\key_mem_ctrl.num_rounds[2] ), .B(\key_reg[3] [16]), 
         .C(n21_adj_8249), .D(n33860), .Z(prev_key0_new_127__N_4659[16])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(85[17:29])
    defparam i1_4_lut_adj_502.init = 16'ha088;
    LUT4 i1_4_lut_adj_503 (.A(\key_mem_ctrl.num_rounds[2] ), .B(\key_reg[3] [17]), 
         .C(n21_adj_8250), .D(n33860), .Z(prev_key0_new_127__N_4659[17])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(85[17:29])
    defparam i1_4_lut_adj_503.init = 16'ha088;
    LUT4 i1_4_lut_adj_504 (.A(\key_mem_ctrl.num_rounds[2] ), .B(\key_reg[3] [18]), 
         .C(n21_adj_8251), .D(n33860), .Z(prev_key0_new_127__N_4659[18])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(85[17:29])
    defparam i1_4_lut_adj_504.init = 16'ha088;
    LUT4 i1_4_lut_adj_505 (.A(\key_mem_ctrl.num_rounds[2] ), .B(\key_reg[3] [19]), 
         .C(n21_adj_8252), .D(n33860), .Z(prev_key0_new_127__N_4659[19])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(85[17:29])
    defparam i1_4_lut_adj_505.init = 16'ha088;
    LUT4 i1_4_lut_adj_506 (.A(\key_mem_ctrl.num_rounds[2] ), .B(\key_reg[3] [20]), 
         .C(n21_adj_8253), .D(n33860), .Z(prev_key0_new_127__N_4659[20])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(85[17:29])
    defparam i1_4_lut_adj_506.init = 16'ha088;
    LUT4 i1_4_lut_adj_507 (.A(\key_mem_ctrl.num_rounds[2] ), .B(\key_reg[3] [21]), 
         .C(n21_adj_8254), .D(n33860), .Z(prev_key0_new_127__N_4659[21])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(85[17:29])
    defparam i1_4_lut_adj_507.init = 16'ha088;
    LUT4 i1_4_lut_adj_508 (.A(\key_mem_ctrl.num_rounds[2] ), .B(\key_reg[3] [22]), 
         .C(n21_adj_8255), .D(n33860), .Z(prev_key0_new_127__N_4659[22])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(85[17:29])
    defparam i1_4_lut_adj_508.init = 16'ha088;
    LUT4 i1_4_lut_adj_509 (.A(\key_mem_ctrl.num_rounds[2] ), .B(\key_reg[3] [23]), 
         .C(n21_adj_8256), .D(n33860), .Z(prev_key0_new_127__N_4659[23])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(85[17:29])
    defparam i1_4_lut_adj_509.init = 16'ha088;
    LUT4 i1_4_lut_adj_510 (.A(\key_mem_ctrl.num_rounds[2] ), .B(\key_reg[3] [24]), 
         .C(n21_adj_8257), .D(n33860), .Z(prev_key0_new_127__N_4659[24])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(85[17:29])
    defparam i1_4_lut_adj_510.init = 16'ha088;
    LUT4 i1_4_lut_adj_511 (.A(\key_mem_ctrl.num_rounds[2] ), .B(\key_reg[3] [25]), 
         .C(n21_adj_8258), .D(n33860), .Z(prev_key0_new_127__N_4659[25])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(85[17:29])
    defparam i1_4_lut_adj_511.init = 16'ha088;
    LUT4 i1_4_lut_adj_512 (.A(\key_mem_ctrl.num_rounds[2] ), .B(\key_reg[3] [26]), 
         .C(n21_adj_8259), .D(n33860), .Z(prev_key0_new_127__N_4659[26])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(85[17:29])
    defparam i1_4_lut_adj_512.init = 16'ha088;
    LUT4 i1_4_lut_adj_513 (.A(\key_mem_ctrl.num_rounds[2] ), .B(\key_reg[3] [27]), 
         .C(n21_adj_8260), .D(n33860), .Z(prev_key0_new_127__N_4659[27])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(85[17:29])
    defparam i1_4_lut_adj_513.init = 16'ha088;
    LUT4 i1_4_lut_adj_514 (.A(\key_mem_ctrl.num_rounds[2] ), .B(\key_reg[3] [28]), 
         .C(n21_adj_8261), .D(n33860), .Z(prev_key0_new_127__N_4659[28])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(85[17:29])
    defparam i1_4_lut_adj_514.init = 16'ha088;
    LUT4 i1_4_lut_adj_515 (.A(\key_mem_ctrl.num_rounds[2] ), .B(\key_reg[3] [29]), 
         .C(n21_adj_8262), .D(n33860), .Z(prev_key0_new_127__N_4659[29])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(85[17:29])
    defparam i1_4_lut_adj_515.init = 16'ha088;
    LUT4 i1_4_lut_adj_516 (.A(\key_mem_ctrl.num_rounds[2] ), .B(\key_reg[3] [30]), 
         .C(n21_adj_8263), .D(n33860), .Z(prev_key0_new_127__N_4659[30])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(85[17:29])
    defparam i1_4_lut_adj_516.init = 16'ha088;
    LUT4 i1_4_lut_adj_517 (.A(\key_mem_ctrl.num_rounds[2] ), .B(\key_reg[3] [31]), 
         .C(n21_adj_8264), .D(n33860), .Z(prev_key0_new_127__N_4659[31])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(85[17:29])
    defparam i1_4_lut_adj_517.init = 16'ha088;
    LUT4 i14570_4_lut (.A(\key_reg[2] [0]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n22), .D(n33860), .Z(prev_key0_new_127__N_4659[32])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14570_4_lut.init = 16'hc088;
    LUT4 i14571_4_lut (.A(\key_reg[2] [1]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n22_adj_8265), .D(n33860), .Z(prev_key0_new_127__N_4659[33])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14571_4_lut.init = 16'hc088;
    LUT4 i14572_4_lut (.A(\key_reg[2] [2]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n22_adj_8266), .D(n33860), .Z(prev_key0_new_127__N_4659[34])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14572_4_lut.init = 16'hc088;
    LUT4 i14573_4_lut (.A(\key_reg[2] [3]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n22_adj_8267), .D(n33860), .Z(prev_key0_new_127__N_4659[35])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14573_4_lut.init = 16'hc088;
    LUT4 i14574_4_lut (.A(\key_reg[2] [4]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n22_adj_8268), .D(n33860), .Z(prev_key0_new_127__N_4659[36])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14574_4_lut.init = 16'hc088;
    LUT4 i14575_4_lut (.A(\key_reg[2] [5]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n22_adj_8269), .D(n33860), .Z(prev_key0_new_127__N_4659[37])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14575_4_lut.init = 16'hc088;
    LUT4 i14576_4_lut (.A(\key_reg[2] [6]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n22_adj_8270), .D(n33860), .Z(prev_key0_new_127__N_4659[38])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14576_4_lut.init = 16'hc088;
    LUT4 i14577_4_lut (.A(\key_reg[2] [7]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n22_adj_8271), .D(n33860), .Z(prev_key0_new_127__N_4659[39])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14577_4_lut.init = 16'hc088;
    LUT4 i14578_4_lut (.A(\key_reg[2] [8]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n22_adj_8272), .D(n33860), .Z(prev_key0_new_127__N_4659[40])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14578_4_lut.init = 16'hc088;
    LUT4 i14579_4_lut (.A(\key_reg[2] [9]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n22_adj_8273), .D(n33860), .Z(prev_key0_new_127__N_4659[41])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14579_4_lut.init = 16'hc088;
    LUT4 i14580_4_lut (.A(\key_reg[2] [10]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n22_adj_8274), .D(n33860), .Z(prev_key0_new_127__N_4659[42])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14580_4_lut.init = 16'hc088;
    LUT4 i14581_4_lut (.A(\key_reg[2] [11]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n22_adj_8275), .D(n33860), .Z(prev_key0_new_127__N_4659[43])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14581_4_lut.init = 16'hc088;
    LUT4 i14582_4_lut (.A(\key_reg[2] [12]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n22_adj_8276), .D(n33860), .Z(prev_key0_new_127__N_4659[44])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14582_4_lut.init = 16'hc088;
    LUT4 i14583_4_lut (.A(\key_reg[2] [13]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n22_adj_8277), .D(n33860), .Z(prev_key0_new_127__N_4659[45])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14583_4_lut.init = 16'hc088;
    LUT4 i14584_4_lut (.A(\key_reg[2] [14]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n22_adj_8278), .D(n33860), .Z(prev_key0_new_127__N_4659[46])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14584_4_lut.init = 16'hc088;
    LUT4 i14585_4_lut (.A(\key_reg[2] [15]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n22_adj_8279), .D(n33860), .Z(prev_key0_new_127__N_4659[47])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14585_4_lut.init = 16'hc088;
    LUT4 i14586_4_lut (.A(\key_reg[2] [16]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n22_adj_8280), .D(n33860), .Z(prev_key0_new_127__N_4659[48])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14586_4_lut.init = 16'hc088;
    LUT4 i14587_4_lut (.A(\key_reg[2] [17]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n22_adj_8281), .D(n33860), .Z(prev_key0_new_127__N_4659[49])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14587_4_lut.init = 16'hc088;
    LUT4 i14588_4_lut (.A(\key_reg[2] [18]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n22_adj_8282), .D(n33860), .Z(prev_key0_new_127__N_4659[50])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14588_4_lut.init = 16'hc088;
    LUT4 i14589_4_lut (.A(\key_reg[2] [19]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n22_adj_8283), .D(n33860), .Z(prev_key0_new_127__N_4659[51])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14589_4_lut.init = 16'hc088;
    LUT4 i14590_4_lut (.A(\key_reg[2] [20]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n22_adj_8284), .D(n33860), .Z(prev_key0_new_127__N_4659[52])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14590_4_lut.init = 16'hc088;
    LUT4 i14591_4_lut (.A(\key_reg[2] [21]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n22_adj_8285), .D(n33860), .Z(prev_key0_new_127__N_4659[53])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14591_4_lut.init = 16'hc088;
    LUT4 i14592_4_lut (.A(\key_reg[2] [22]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n22_adj_8286), .D(n33860), .Z(prev_key0_new_127__N_4659[54])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14592_4_lut.init = 16'hc088;
    LUT4 i14593_4_lut (.A(\key_reg[2] [23]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n22_adj_8287), .D(n33860), .Z(prev_key0_new_127__N_4659[55])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14593_4_lut.init = 16'hc088;
    LUT4 i14594_4_lut (.A(\key_reg[2] [24]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n22_adj_8288), .D(n33860), .Z(prev_key0_new_127__N_4659[56])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14594_4_lut.init = 16'hc088;
    LUT4 i14595_4_lut (.A(\key_reg[2] [25]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n22_adj_8289), .D(n33860), .Z(prev_key0_new_127__N_4659[57])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14595_4_lut.init = 16'hc088;
    LUT4 i14596_4_lut (.A(\key_reg[2] [26]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n22_adj_8290), .D(n33860), .Z(prev_key0_new_127__N_4659[58])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14596_4_lut.init = 16'hc088;
    LUT4 i14597_4_lut (.A(\key_reg[2] [27]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n22_adj_8291), .D(n33860), .Z(prev_key0_new_127__N_4659[59])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14597_4_lut.init = 16'hc088;
    LUT4 i1_3_lut_4_lut_rep_694 (.A(n33943), .B(n33944), .C(\key_mem_ctrl.num_rounds[2] ), 
         .D(n28850), .Z(clk_c_enable_2335)) /* synthesis lut_function=(A (D)+!A (B (D)+!B !(C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_3_lut_4_lut_rep_694.init = 16'hef00;
    LUT4 i14598_4_lut (.A(\key_reg[2] [28]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n22_adj_8292), .D(n33860), .Z(prev_key0_new_127__N_4659[60])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14598_4_lut.init = 16'hc088;
    LUT4 i14599_4_lut (.A(\key_reg[2] [29]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n22_adj_8293), .D(n33860), .Z(prev_key0_new_127__N_4659[61])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14599_4_lut.init = 16'hc088;
    LUT4 i14600_4_lut (.A(\key_reg[2] [30]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n22_adj_8294), .D(n33860), .Z(prev_key0_new_127__N_4659[62])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14600_4_lut.init = 16'hc088;
    LUT4 i14601_4_lut (.A(\key_reg[2] [31]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n22_adj_8295), .D(n33860), .Z(prev_key0_new_127__N_4659[63])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14601_4_lut.init = 16'hc088;
    LUT4 i14602_4_lut (.A(\key_reg[1] [0]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[64]), .D(n33860), .Z(prev_key0_new_127__N_4659[64])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14602_4_lut.init = 16'hc088;
    LUT4 i14603_4_lut (.A(\key_reg[1] [1]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[65]), .D(n33860), .Z(prev_key0_new_127__N_4659[65])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14603_4_lut.init = 16'hc088;
    LUT4 i14604_4_lut (.A(\key_reg[1] [2]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[66]), .D(n33860), .Z(prev_key0_new_127__N_4659[66])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14604_4_lut.init = 16'hc088;
    LUT4 i14605_4_lut (.A(\key_reg[1] [3]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[67]), .D(n33860), .Z(prev_key0_new_127__N_4659[67])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14605_4_lut.init = 16'hc088;
    LUT4 i14606_4_lut (.A(\key_reg[1] [4]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[68]), .D(n33860), .Z(prev_key0_new_127__N_4659[68])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14606_4_lut.init = 16'hc088;
    LUT4 i1_3_lut_4_lut_rep_695 (.A(n33943), .B(n33944), .C(\key_mem_ctrl.num_rounds[2] ), 
         .D(n28850), .Z(clk_c_enable_2385)) /* synthesis lut_function=(A (D)+!A (B (D)+!B !(C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_3_lut_4_lut_rep_695.init = 16'hef00;
    LUT4 i14607_4_lut (.A(\key_reg[1] [5]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[69]), .D(n33860), .Z(prev_key0_new_127__N_4659[69])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14607_4_lut.init = 16'hc088;
    LUT4 i14608_4_lut (.A(\key_reg[1] [6]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[70]), .D(n33860), .Z(prev_key0_new_127__N_4659[70])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14608_4_lut.init = 16'hc088;
    LUT4 i14609_4_lut (.A(\key_reg[1] [7]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[71]), .D(n33860), .Z(prev_key0_new_127__N_4659[71])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14609_4_lut.init = 16'hc088;
    LUT4 i14610_4_lut (.A(\key_reg[1] [8]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[72]), .D(n33860), .Z(prev_key0_new_127__N_4659[72])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14610_4_lut.init = 16'hc088;
    LUT4 i14611_4_lut (.A(\key_reg[1] [9]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[73]), .D(n33860), .Z(prev_key0_new_127__N_4659[73])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14611_4_lut.init = 16'hc088;
    LUT4 i14612_4_lut (.A(\key_reg[1] [10]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[74]), .D(n33860), .Z(prev_key0_new_127__N_4659[74])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14612_4_lut.init = 16'hc088;
    LUT4 i14613_4_lut (.A(\key_reg[1] [11]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[75]), .D(n33860), .Z(prev_key0_new_127__N_4659[75])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14613_4_lut.init = 16'hc088;
    LUT4 i14614_4_lut (.A(\key_reg[1] [12]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[76]), .D(n33860), .Z(prev_key0_new_127__N_4659[76])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14614_4_lut.init = 16'hc088;
    LUT4 i14615_4_lut (.A(\key_reg[1] [13]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[77]), .D(n33860), .Z(prev_key0_new_127__N_4659[77])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14615_4_lut.init = 16'hc088;
    LUT4 i14616_4_lut (.A(\key_reg[1] [14]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[78]), .D(n33860), .Z(prev_key0_new_127__N_4659[78])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14616_4_lut.init = 16'hc088;
    LUT4 i14617_4_lut (.A(\key_reg[1] [15]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[79]), .D(n33860), .Z(prev_key0_new_127__N_4659[79])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14617_4_lut.init = 16'hc088;
    LUT4 i14618_4_lut (.A(\key_reg[1] [16]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[80]), .D(n33860), .Z(prev_key0_new_127__N_4659[80])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14618_4_lut.init = 16'hc088;
    LUT4 i14619_4_lut (.A(\key_reg[1] [17]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[81]), .D(n33860), .Z(prev_key0_new_127__N_4659[81])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14619_4_lut.init = 16'hc088;
    LUT4 i14620_4_lut (.A(\key_reg[1] [18]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[82]), .D(n33860), .Z(prev_key0_new_127__N_4659[82])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14620_4_lut.init = 16'hc088;
    LUT4 i14621_4_lut (.A(\key_reg[1] [19]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[83]), .D(n33860), .Z(prev_key0_new_127__N_4659[83])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14621_4_lut.init = 16'hc088;
    LUT4 i14622_4_lut (.A(\key_reg[1] [20]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[84]), .D(n33860), .Z(prev_key0_new_127__N_4659[84])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14622_4_lut.init = 16'hc088;
    LUT4 round_3__I_0_Mux_98_i11_3_lut (.A(\key_mem[12] [98]), .B(\key_mem[13] [98]), 
         .C(n33952), .Z(n11_adj_1)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_98_i11_3_lut.init = 16'hcaca;
    LUT4 i14623_4_lut (.A(\key_reg[1] [21]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[85]), .D(n33860), .Z(prev_key0_new_127__N_4659[85])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14623_4_lut.init = 16'hc088;
    LUT4 i14624_4_lut (.A(\key_reg[1] [22]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[86]), .D(n33860), .Z(prev_key0_new_127__N_4659[86])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14624_4_lut.init = 16'hc088;
    LUT4 round_3__I_0_Mux_98_i9_3_lut (.A(\key_mem[10] [98]), .B(\key_mem[11] [98]), 
         .C(n33952), .Z(n9_adj_8308)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_98_i9_3_lut.init = 16'hcaca;
    LUT4 i14625_4_lut (.A(\key_reg[1] [23]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[87]), .D(n33860), .Z(prev_key0_new_127__N_4659[87])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14625_4_lut.init = 16'hc088;
    LUT4 i14626_4_lut (.A(\key_reg[1] [24]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[88]), .D(n33860), .Z(prev_key0_new_127__N_4659[88])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14626_4_lut.init = 16'hc088;
    LUT4 i14627_4_lut (.A(\key_reg[1] [25]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[89]), .D(n33860), .Z(prev_key0_new_127__N_4659[89])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14627_4_lut.init = 16'hc088;
    LUT4 i14628_4_lut (.A(\key_reg[1] [26]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[90]), .D(n33860), .Z(prev_key0_new_127__N_4659[90])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14628_4_lut.init = 16'hc088;
    LUT4 i14629_4_lut (.A(\key_reg[1] [27]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[91]), .D(n33860), .Z(prev_key0_new_127__N_4659[91])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14629_4_lut.init = 16'hc088;
    LUT4 i14630_4_lut (.A(\key_reg[1] [28]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[92]), .D(n33860), .Z(prev_key0_new_127__N_4659[92])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14630_4_lut.init = 16'hc088;
    LUT4 i14631_4_lut (.A(\key_reg[1] [29]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[93]), .D(n33860), .Z(prev_key0_new_127__N_4659[93])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14631_4_lut.init = 16'hc088;
    LUT4 i14632_4_lut (.A(\key_reg[1] [30]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[94]), .D(n33860), .Z(prev_key0_new_127__N_4659[94])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14632_4_lut.init = 16'hc088;
    LUT4 i14633_4_lut (.A(\key_reg[1] [31]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[95]), .D(n33860), .Z(prev_key0_new_127__N_4659[95])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14633_4_lut.init = 16'hc088;
    LUT4 new_sboxw_23__I_0_i30_2_lut_rep_414 (.A(\new_sboxw[21] ), .B(\rcon_logic.tmp_rcon [6]), 
         .Z(n33718)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(224[13:27])
    defparam new_sboxw_23__I_0_i30_2_lut_rep_414.init = 16'h6666;
    LUT4 i14634_4_lut (.A(\key_reg[0] [0]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[96]), .D(n33860), .Z(prev_key0_new_127__N_4659[96])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14634_4_lut.init = 16'hc088;
    LUT4 i14635_4_lut (.A(\key_reg[0] [1]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[97]), .D(n33860), .Z(prev_key0_new_127__N_4659[97])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14635_4_lut.init = 16'hc088;
    LUT4 i14636_4_lut (.A(\key_reg[0] [2]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[98]), .D(n33860), .Z(prev_key0_new_127__N_4659[98])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14636_4_lut.init = 16'hc088;
    LUT4 i14637_4_lut (.A(\key_reg[0] [3]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[99]), .D(n33860), .Z(prev_key0_new_127__N_4659[99])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14637_4_lut.init = 16'hc088;
    LUT4 i14638_4_lut (.A(\key_reg[0] [4]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[100]), .D(n33860), .Z(prev_key0_new_127__N_4659[100])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14638_4_lut.init = 16'hc088;
    LUT4 i14639_4_lut (.A(\key_reg[0] [5]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[101]), .D(n33860), .Z(prev_key0_new_127__N_4659[101])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14639_4_lut.init = 16'hc088;
    LUT4 mux_85_i75_3_lut_rep_243_4_lut (.A(prev_key0_reg[74]), .B(n4), 
         .C(n33859), .D(\key_reg[5] [10]), .Z(n33547)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam mux_85_i75_3_lut_rep_243_4_lut.init = 16'h6f60;
    LUT4 i14640_4_lut (.A(\key_reg[0] [6]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[102]), .D(n33860), .Z(prev_key0_new_127__N_4659[102])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14640_4_lut.init = 16'hc088;
    LUT4 round_3__I_0_Mux_98_i8_3_lut (.A(\key_mem[8] [98]), .B(\key_mem[9] [98]), 
         .C(n33952), .Z(n8_adj_8315)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_98_i8_3_lut.init = 16'hcaca;
    LUT4 i14641_4_lut (.A(\key_reg[0] [7]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[103]), .D(n33860), .Z(prev_key0_new_127__N_4659[103])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14641_4_lut.init = 16'hc088;
    LUT4 i2_3_lut_rep_311_4_lut (.A(\new_sboxw[21] ), .B(\rcon_logic.tmp_rcon [6]), 
         .C(prev_key1_reg[125]), .D(prev_key1_reg[93]), .Z(n33615)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(224[13:27])
    defparam i2_3_lut_rep_311_4_lut.init = 16'h6996;
    LUT4 round_3__I_0_Mux_98_i5_3_lut (.A(\key_mem[6] [98]), .B(\key_mem[7] [98]), 
         .C(n33952), .Z(n5_adj_8316)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_98_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_98_i4_3_lut (.A(\key_mem[4] [98]), .B(\key_mem[5] [98]), 
         .C(n33952), .Z(n4_adj_8317)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_98_i4_3_lut.init = 16'hcaca;
    LUT4 i14642_4_lut (.A(\key_reg[0] [8]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[104]), .D(n33860), .Z(prev_key0_new_127__N_4659[104])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14642_4_lut.init = 16'hc088;
    LUT4 new_sboxw_23__I_0_i29_2_lut_rep_415 (.A(\new_sboxw[20] ), .B(\rcon_logic.tmp_rcon [5]), 
         .Z(n33719)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(224[13:27])
    defparam new_sboxw_23__I_0_i29_2_lut_rep_415.init = 16'h6666;
    LUT4 i14643_4_lut (.A(\key_reg[0] [9]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[105]), .D(n33860), .Z(prev_key0_new_127__N_4659[105])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14643_4_lut.init = 16'hc088;
    LUT4 i14644_4_lut (.A(\key_reg[0] [10]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[106]), .D(n33860), .Z(prev_key0_new_127__N_4659[106])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14644_4_lut.init = 16'hc088;
    LUT4 i14645_4_lut (.A(\key_reg[0] [11]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[107]), .D(n33860), .Z(prev_key0_new_127__N_4659[107])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14645_4_lut.init = 16'hc088;
    LUT4 i14646_4_lut (.A(\key_reg[0] [12]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[108]), .D(n33860), .Z(prev_key0_new_127__N_4659[108])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14646_4_lut.init = 16'hc088;
    LUT4 i14647_4_lut (.A(\key_reg[0] [13]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[109]), .D(n33860), .Z(prev_key0_new_127__N_4659[109])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14647_4_lut.init = 16'hc088;
    LUT4 i14648_4_lut (.A(\key_reg[0] [14]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[110]), .D(n33860), .Z(prev_key0_new_127__N_4659[110])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14648_4_lut.init = 16'hc088;
    LUT4 i14649_4_lut (.A(\key_reg[0] [15]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[111]), .D(n33860), .Z(prev_key0_new_127__N_4659[111])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14649_4_lut.init = 16'hc088;
    LUT4 i14650_4_lut (.A(\key_reg[0] [16]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[112]), .D(n33860), .Z(prev_key0_new_127__N_4659[112])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14650_4_lut.init = 16'hc088;
    LUT4 i14651_4_lut (.A(\key_reg[0] [17]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[113]), .D(n33860), .Z(prev_key0_new_127__N_4659[113])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14651_4_lut.init = 16'hc088;
    LUT4 i14652_4_lut (.A(\key_reg[0] [18]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[114]), .D(n33860), .Z(prev_key0_new_127__N_4659[114])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14652_4_lut.init = 16'hc088;
    LUT4 i14653_4_lut (.A(\key_reg[0] [19]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[115]), .D(n33860), .Z(prev_key0_new_127__N_4659[115])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14653_4_lut.init = 16'hc088;
    LUT4 i14654_4_lut (.A(\key_reg[0] [20]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[116]), .D(n33860), .Z(prev_key0_new_127__N_4659[116])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14654_4_lut.init = 16'hc088;
    LUT4 i14655_4_lut (.A(\key_reg[0] [21]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[117]), .D(n33860), .Z(prev_key0_new_127__N_4659[117])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14655_4_lut.init = 16'hc088;
    LUT4 i14656_4_lut (.A(\key_reg[0] [22]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[118]), .D(n33860), .Z(prev_key0_new_127__N_4659[118])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14656_4_lut.init = 16'hc088;
    LUT4 i14657_4_lut (.A(\key_reg[0] [23]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[119]), .D(n33860), .Z(prev_key0_new_127__N_4659[119])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14657_4_lut.init = 16'hc088;
    LUT4 i14658_4_lut (.A(\key_reg[0] [24]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[120]), .D(n33860), .Z(prev_key0_new_127__N_4659[120])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14658_4_lut.init = 16'hc088;
    LUT4 i2_3_lut_rep_312_4_lut (.A(\new_sboxw[20] ), .B(\rcon_logic.tmp_rcon [5]), 
         .C(prev_key1_reg[124]), .D(prev_key1_reg[92]), .Z(n33616)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(224[13:27])
    defparam i2_3_lut_rep_312_4_lut.init = 16'h6996;
    LUT4 i14659_4_lut (.A(\key_reg[0] [25]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[121]), .D(n33860), .Z(prev_key0_new_127__N_4659[121])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14659_4_lut.init = 16'hc088;
    LUT4 i14660_4_lut (.A(\key_reg[0] [26]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[122]), .D(n33860), .Z(prev_key0_new_127__N_4659[122])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14660_4_lut.init = 16'hc088;
    LUT4 i14661_4_lut (.A(\key_reg[0] [27]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[123]), .D(n33860), .Z(prev_key0_new_127__N_4659[123])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14661_4_lut.init = 16'hc088;
    LUT4 i14662_4_lut (.A(\key_reg[0] [28]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[124]), .D(n33860), .Z(prev_key0_new_127__N_4659[124])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14662_4_lut.init = 16'hc088;
    LUT4 i14663_4_lut (.A(\key_reg[0] [29]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[125]), .D(n33860), .Z(prev_key0_new_127__N_4659[125])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14663_4_lut.init = 16'hc088;
    LUT4 i14664_4_lut (.A(\key_reg[0] [30]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[126]), .D(n33860), .Z(prev_key0_new_127__N_4659[126])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14664_4_lut.init = 16'hc088;
    LUT4 i14665_4_lut (.A(\key_reg[0] [31]), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n8680[127]), .D(n33860), .Z(prev_key0_new_127__N_4659[127])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i14665_4_lut.init = 16'hc088;
    LUT4 i6_2_lut_3_lut (.A(prev_key1_reg[41]), .B(n33738), .C(keymem_sboxw[9]), 
         .Z(n15897)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;
    defparam i6_2_lut_3_lut.init = 16'h9696;
    LUT4 i1_3_lut (.A(n35839), .B(\rcon_logic.tmp_rcon [2]), .C(n72), 
         .Z(rcon_new[2])) /* synthesis lut_function=((B (C))+!A) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam i1_3_lut.init = 16'hd5d5;
    LUT4 i1_4_lut_adj_518 (.A(n35839), .B(rcon_reg[2]), .C(n72), .D(\rcon_logic.tmp_rcon [0]), 
         .Z(rcon_new[3])) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam i1_4_lut_adj_518.init = 16'h75d5;
    LUT4 i1_3_lut_adj_519 (.A(n35839), .B(\rcon_logic.tmp_rcon [7]), .C(n72), 
         .Z(rcon_new[7])) /* synthesis lut_function=((B (C))+!A) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam i1_3_lut_adj_519.init = 16'hd5d5;
    LUT4 round_3__I_0_Mux_98_i2_3_lut (.A(\key_mem[2] [98]), .B(\key_mem[3] [98]), 
         .C(n33952), .Z(n2_adj_8318)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_98_i2_3_lut.init = 16'hcaca;
    LUT4 i6_2_lut_3_lut_adj_520 (.A(prev_key1_reg[32]), .B(n33747), .C(keymem_sboxw[0]), 
         .Z(n15304)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;
    defparam i6_2_lut_3_lut_adj_520.init = 16'h9696;
    LUT4 new_sboxw_23__I_0_i28_2_lut_rep_416 (.A(\new_sboxw[19] ), .B(rcon_reg[3]), 
         .Z(n33720)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(224[13:27])
    defparam new_sboxw_23__I_0_i28_2_lut_rep_416.init = 16'h6666;
    LUT4 round_3__I_0_Mux_98_i1_3_lut (.A(\key_mem[0] [98]), .B(\key_mem[1] [98]), 
         .C(n33952), .Z(n1_adj_8319)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_98_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_115_i11_3_lut (.A(\key_mem[12] [115]), .B(\key_mem[13] [115]), 
         .C(n33952), .Z(n11_adj_2)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_115_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_115_i9_3_lut (.A(\key_mem[10] [115]), .B(\key_mem[11] [115]), 
         .C(n33952), .Z(n9_adj_8321)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_115_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_115_i8_3_lut (.A(\key_mem[8] [115]), .B(\key_mem[9] [115]), 
         .C(n33952), .Z(n8_adj_8322)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_115_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_115_i5_3_lut (.A(\key_mem[6] [115]), .B(\key_mem[7] [115]), 
         .C(n33952), .Z(n5_adj_8323)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_115_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_115_i4_3_lut (.A(\key_mem[4] [115]), .B(\key_mem[5] [115]), 
         .C(n33952), .Z(n4_adj_8324)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_115_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_115_i2_3_lut (.A(\key_mem[2] [115]), .B(\key_mem[3] [115]), 
         .C(n33952), .Z(n2_adj_8325)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_115_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_115_i1_3_lut (.A(\key_mem[0] [115]), .B(\key_mem[1] [115]), 
         .C(n33952), .Z(n1_adj_8326)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_115_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_114_i11_3_lut (.A(\key_mem[12] [114]), .B(\key_mem[13] [114]), 
         .C(n33952), .Z(n11_adj_3)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_114_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_88_i2_3_lut (.A(\key_mem[2] [88]), .B(\key_mem[3] [88]), 
         .C(n33952), .Z(n2_adj_8328)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_88_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_114_i9_3_lut (.A(\key_mem[10] [114]), .B(\key_mem[11] [114]), 
         .C(n33952), .Z(n9_adj_8329)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_114_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_114_i8_3_lut (.A(\key_mem[8] [114]), .B(\key_mem[9] [114]), 
         .C(n33952), .Z(n8_adj_8330)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_114_i8_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_521 (.A(n33860), .B(n33667), .C(n15314), .D(n35835), 
         .Z(n15316)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_4_lut_adj_521.init = 16'ha088;
    LUT4 i9706_4_lut (.A(\key_reg[6] [0]), .B(prev_key0_reg[32]), .C(n33859), 
         .D(n33666), .Z(n15314)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i9706_4_lut.init = 16'h3aca;
    LUT4 i3049_4_lut (.A(prev_key0_reg[96]), .B(\round_key_gen.trw[0] ), 
         .C(\round_key_gen.trw[8] ), .D(n35834), .Z(n8487)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)))+!A !(B (C+!(D))+!B (C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i3049_4_lut.init = 16'h5a66;
    LUT4 round_3__I_0_Mux_88_i1_3_lut (.A(\key_mem[0] [88]), .B(\key_mem[1] [88]), 
         .C(n33952), .Z(n1_adj_8331)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_88_i1_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_522 (.A(n33860), .B(n33664), .C(n15427), .D(n35835), 
         .Z(n15429)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_4_lut_adj_522.init = 16'ha088;
    LUT4 i9821_4_lut (.A(\key_reg[6] [1]), .B(prev_key0_reg[33]), .C(n33859), 
         .D(n33665), .Z(n15427)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i9821_4_lut.init = 16'h3aca;
    LUT4 i3443_4_lut (.A(prev_key0_reg[97]), .B(\round_key_gen.trw[1] ), 
         .C(\round_key_gen.trw[9] ), .D(n35834), .Z(n8929)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)))+!A !(B (C+!(D))+!B (C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i3443_4_lut.init = 16'h5a66;
    LUT4 i1_4_lut_adj_523 (.A(n33860), .B(n33662), .C(n15487), .D(n35835), 
         .Z(n15489)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_4_lut_adj_523.init = 16'ha088;
    LUT4 i9882_4_lut (.A(\key_reg[6] [2]), .B(prev_key0_reg[34]), .C(n33859), 
         .D(n33663), .Z(n15487)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i9882_4_lut.init = 16'h3aca;
    LUT4 i1_4_lut_adj_524 (.A(prev_key0_reg[98]), .B(\round_key_gen.trw[2] ), 
         .C(\round_key_gen.trw[10] ), .D(n35834), .Z(n4_adj_8332)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)))+!A !(B (C+!(D))+!B (C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i1_4_lut_adj_524.init = 16'h5a66;
    LUT4 i1_4_lut_adj_525 (.A(n33860), .B(n33660), .C(n15547), .D(n35835), 
         .Z(n15549)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_4_lut_adj_525.init = 16'ha088;
    LUT4 i9943_4_lut (.A(\key_reg[6] [3]), .B(prev_key0_reg[35]), .C(n33859), 
         .D(n33661), .Z(n15547)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i9943_4_lut.init = 16'h3aca;
    LUT4 i1_4_lut_adj_526 (.A(prev_key0_reg[99]), .B(\round_key_gen.trw[3] ), 
         .C(\round_key_gen.trw[11] ), .D(n35834), .Z(n4_adj_8333)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)))+!A !(B (C+!(D))+!B (C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i1_4_lut_adj_526.init = 16'h5a66;
    LUT4 i1_4_lut_adj_527 (.A(n33860), .B(n33658), .C(n15607), .D(n35835), 
         .Z(n15609)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_4_lut_adj_527.init = 16'ha088;
    LUT4 i10004_4_lut (.A(\key_reg[6] [4]), .B(prev_key0_reg[36]), .C(n33859), 
         .D(n33659), .Z(n15607)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i10004_4_lut.init = 16'h3aca;
    LUT4 round_3__I_0_Mux_87_i11_3_lut (.A(\key_mem[12] [87]), .B(\key_mem[13] [87]), 
         .C(n33952), .Z(n11_adj_4)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_87_i11_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_528 (.A(prev_key0_reg[100]), .B(\round_key_gen.trw[4] ), 
         .C(\round_key_gen.trw[12] ), .D(n35834), .Z(n4_adj_8335)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)))+!A !(B (C+!(D))+!B (C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i1_4_lut_adj_528.init = 16'h5a66;
    LUT4 i1_4_lut_adj_529 (.A(n33860), .B(n33656), .C(n15667), .D(n35835), 
         .Z(n15669)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_4_lut_adj_529.init = 16'ha088;
    LUT4 i10065_4_lut (.A(\key_reg[6] [5]), .B(prev_key0_reg[37]), .C(n33859), 
         .D(n33657), .Z(n15667)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i10065_4_lut.init = 16'h3aca;
    LUT4 i1_4_lut_adj_530 (.A(prev_key0_reg[101]), .B(\round_key_gen.trw[5] ), 
         .C(\round_key_gen.trw[13] ), .D(n35834), .Z(n4_adj_8336)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)))+!A !(B (C+!(D))+!B (C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i1_4_lut_adj_530.init = 16'h5a66;
    LUT4 i1_4_lut_adj_531 (.A(n33860), .B(n33654), .C(n15727), .D(n35835), 
         .Z(n15729)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_4_lut_adj_531.init = 16'ha088;
    LUT4 i10126_4_lut (.A(\key_reg[6] [6]), .B(prev_key0_reg[38]), .C(n33859), 
         .D(n33655), .Z(n15727)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i10126_4_lut.init = 16'h3aca;
    LUT4 i1_4_lut_adj_532 (.A(prev_key0_reg[102]), .B(\round_key_gen.trw[6] ), 
         .C(\round_key_gen.trw[14] ), .D(n35834), .Z(n4_adj_8337)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)))+!A !(B (C+!(D))+!B (C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i1_4_lut_adj_532.init = 16'h5a66;
    LUT4 i1_4_lut_adj_533 (.A(n33860), .B(n33652), .C(n15787), .D(n35835), 
         .Z(n15789)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_4_lut_adj_533.init = 16'ha088;
    LUT4 i10187_4_lut (.A(\key_reg[6] [7]), .B(prev_key0_reg[39]), .C(n33859), 
         .D(n33653), .Z(n15787)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i10187_4_lut.init = 16'h3aca;
    LUT4 round_3__I_0_Mux_87_i9_3_lut (.A(\key_mem[10] [87]), .B(\key_mem[11] [87]), 
         .C(n33952), .Z(n9_adj_8338)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_87_i9_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_534 (.A(prev_key0_reg[103]), .B(\round_key_gen.trw[7] ), 
         .C(\round_key_gen.trw[15] ), .D(n35834), .Z(n4_adj_8339)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)))+!A !(B (C+!(D))+!B (C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i1_4_lut_adj_534.init = 16'h5a66;
    LUT4 round_3__I_0_Mux_87_i8_3_lut (.A(\key_mem[8] [87]), .B(\key_mem[9] [87]), 
         .C(n33952), .Z(n8_adj_8340)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_87_i8_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_rep_313_4_lut (.A(\new_sboxw[19] ), .B(rcon_reg[3]), .C(prev_key1_reg[123]), 
         .D(prev_key1_reg[91]), .Z(n33617)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(224[13:27])
    defparam i2_3_lut_rep_313_4_lut.init = 16'h6996;
    LUT4 i1_4_lut_adj_535 (.A(n33860), .B(n33650), .C(n15847), .D(n35835), 
         .Z(n15849)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_4_lut_adj_535.init = 16'ha088;
    LUT4 i10248_4_lut (.A(\key_reg[6] [8]), .B(prev_key0_reg[40]), .C(n33859), 
         .D(n33651), .Z(n15847)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i10248_4_lut.init = 16'h3aca;
    LUT4 round_3__I_0_Mux_114_i5_3_lut (.A(\key_mem[6] [114]), .B(\key_mem[7] [114]), 
         .C(n33952), .Z(n5_adj_8341)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_114_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_114_i4_3_lut (.A(\key_mem[4] [114]), .B(\key_mem[5] [114]), 
         .C(n33952), .Z(n4_adj_8342)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_114_i4_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_536 (.A(prev_key0_reg[104]), .B(\round_key_gen.trw[8] ), 
         .C(\round_key_gen.trw[16] ), .D(n35834), .Z(n4_adj_8343)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)))+!A !(B (C+!(D))+!B (C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i1_4_lut_adj_536.init = 16'h5a66;
    LUT4 round_3__I_0_Mux_114_i2_3_lut (.A(\key_mem[2] [114]), .B(\key_mem[3] [114]), 
         .C(n33952), .Z(n2_adj_8344)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_114_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_114_i1_3_lut (.A(\key_mem[0] [114]), .B(\key_mem[1] [114]), 
         .C(n33952), .Z(n1_adj_8345)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_114_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_97_i11_3_lut (.A(\key_mem[12] [97]), .B(\key_mem[13] [97]), 
         .C(n33952), .Z(n11_adj_5)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_97_i11_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_537 (.A(n33860), .B(n33648), .C(n15907), .D(n35835), 
         .Z(n15909)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_4_lut_adj_537.init = 16'ha088;
    LUT4 i10309_4_lut (.A(\key_reg[6] [9]), .B(prev_key0_reg[41]), .C(n33859), 
         .D(n33649), .Z(n15907)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i10309_4_lut.init = 16'h3aca;
    LUT4 round_3__I_0_Mux_113_i11_3_lut (.A(\key_mem[12] [113]), .B(\key_mem[13] [113]), 
         .C(n33952), .Z(n11_adj_6)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_113_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_97_i9_3_lut (.A(\key_mem[10] [97]), .B(\key_mem[11] [97]), 
         .C(n33952), .Z(n9_adj_8348)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_97_i9_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_538 (.A(prev_key0_reg[105]), .B(\round_key_gen.trw[9] ), 
         .C(\round_key_gen.trw[17] ), .D(n35834), .Z(n4_adj_8349)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)))+!A !(B (C+!(D))+!B (C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i1_4_lut_adj_538.init = 16'h5a66;
    LUT4 round_3__I_0_Mux_97_i8_3_lut (.A(\key_mem[8] [97]), .B(\key_mem[9] [97]), 
         .C(n33952), .Z(n8_adj_8350)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_97_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_87_i5_3_lut (.A(\key_mem[6] [87]), .B(\key_mem[7] [87]), 
         .C(n33952), .Z(n5_adj_8351)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_87_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_113_i9_3_lut (.A(\key_mem[10] [113]), .B(\key_mem[11] [113]), 
         .C(n33952), .Z(n9_adj_8352)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_113_i9_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_539 (.A(n33860), .B(n33646), .C(n15967), .D(n35835), 
         .Z(n15969)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_4_lut_adj_539.init = 16'ha088;
    LUT4 round_3__I_0_Mux_113_i8_3_lut (.A(\key_mem[8] [113]), .B(\key_mem[9] [113]), 
         .C(n33952), .Z(n8_adj_8353)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_113_i8_3_lut.init = 16'hcaca;
    LUT4 i10370_4_lut (.A(\key_reg[6] [10]), .B(prev_key0_reg[42]), .C(n33859), 
         .D(n33647), .Z(n15967)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i10370_4_lut.init = 16'h3aca;
    LUT4 round_3__I_0_Mux_87_i4_3_lut (.A(\key_mem[4] [87]), .B(\key_mem[5] [87]), 
         .C(n33952), .Z(n4_adj_8354)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_87_i4_3_lut.init = 16'hcaca;
    LUT4 i2_2_lut_rep_345 (.A(prev_key0_reg[73]), .B(n4_adj_8349), .Z(n33649)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i2_2_lut_rep_345.init = 16'h6666;
    LUT4 round_3__I_0_Mux_113_i5_3_lut (.A(\key_mem[6] [113]), .B(\key_mem[7] [113]), 
         .C(n33952), .Z(n5_adj_8355)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_113_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_97_i5_3_lut (.A(\key_mem[6] [97]), .B(\key_mem[7] [97]), 
         .C(n33952), .Z(n5_adj_8356)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_97_i5_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_540 (.A(prev_key0_reg[106]), .B(\round_key_gen.trw[10] ), 
         .C(\round_key_gen.trw[18] ), .D(n35834), .Z(n4)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)))+!A !(B (C+!(D))+!B (C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i1_4_lut_adj_540.init = 16'h5a66;
    LUT4 round_3__I_0_Mux_113_i4_3_lut (.A(\key_mem[4] [113]), .B(\key_mem[5] [113]), 
         .C(n33952), .Z(n4_adj_8357)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_113_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_113_i2_3_lut (.A(\key_mem[2] [113]), .B(\key_mem[3] [113]), 
         .C(n33952), .Z(n2_adj_8358)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_113_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_97_i4_3_lut (.A(\key_mem[4] [97]), .B(\key_mem[5] [97]), 
         .C(n33952), .Z(n4_adj_8359)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_97_i4_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_541 (.A(n33860), .B(n33644), .C(n16027), .D(n35835), 
         .Z(n16029)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_4_lut_adj_541.init = 16'ha088;
    LUT4 new_sboxw_23__I_0_i27_2_lut_rep_417 (.A(\new_sboxw[18] ), .B(rcon_reg[2]), 
         .Z(n33721)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(224[13:27])
    defparam new_sboxw_23__I_0_i27_2_lut_rep_417.init = 16'h6666;
    LUT4 mux_85_i74_3_lut_rep_244_4_lut (.A(prev_key0_reg[73]), .B(n4_adj_8349), 
         .C(n33859), .D(\key_reg[5] [9]), .Z(n33548)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam mux_85_i74_3_lut_rep_244_4_lut.init = 16'h6f60;
    LUT4 i2_3_lut_rep_314_4_lut (.A(\new_sboxw[18] ), .B(rcon_reg[2]), .C(prev_key1_reg[122]), 
         .D(prev_key1_reg[90]), .Z(n33618)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(224[13:27])
    defparam i2_3_lut_rep_314_4_lut.init = 16'h6996;
    LUT4 i10431_4_lut (.A(\key_reg[6] [11]), .B(prev_key0_reg[43]), .C(n33859), 
         .D(n33645), .Z(n16027)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i10431_4_lut.init = 16'h3aca;
    LUT4 round_3__I_0_Mux_113_i1_3_lut (.A(\key_mem[0] [113]), .B(\key_mem[1] [113]), 
         .C(n33952), .Z(n1_adj_8360)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_113_i1_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_542 (.A(prev_key0_reg[107]), .B(\round_key_gen.trw[11] ), 
         .C(\round_key_gen.trw[19] ), .D(n35834), .Z(n4_adj_8361)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)))+!A !(B (C+!(D))+!B (C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i1_4_lut_adj_542.init = 16'h5a66;
    LUT4 i2_3_lut_rep_418 (.A(\new_sboxw[17] ), .B(prev_key1_reg[121]), 
         .C(\rcon_logic.tmp_rcon [2]), .Z(n33722)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(110[18:27])
    defparam i2_3_lut_rep_418.init = 16'h9696;
    LUT4 round_3__I_0_Mux_87_i2_3_lut (.A(\key_mem[2] [87]), .B(\key_mem[3] [87]), 
         .C(n33952), .Z(n2_adj_8362)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_87_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_112_i11_3_lut (.A(\key_mem[12] [112]), .B(\key_mem[13] [112]), 
         .C(n33952), .Z(n11_adj_7)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_112_i11_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_543 (.A(n33860), .B(n33642), .C(n16087), .D(n35835), 
         .Z(n16089)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_4_lut_adj_543.init = 16'ha088;
    LUT4 round_3__I_0_Mux_112_i9_3_lut (.A(\key_mem[10] [112]), .B(\key_mem[11] [112]), 
         .C(n33952), .Z(n9_adj_8364)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_112_i9_3_lut.init = 16'hcaca;
    LUT4 i10492_4_lut (.A(\key_reg[6] [12]), .B(prev_key0_reg[44]), .C(n33859), 
         .D(n33643), .Z(n16087)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i10492_4_lut.init = 16'h3aca;
    LUT4 round_3__I_0_Mux_97_i2_3_lut (.A(\key_mem[2] [97]), .B(\key_mem[3] [97]), 
         .C(n33952), .Z(n2_adj_8365)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_97_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_112_i8_3_lut (.A(\key_mem[8] [112]), .B(\key_mem[9] [112]), 
         .C(n33952), .Z(n8_adj_8366)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_112_i8_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_544 (.A(prev_key0_reg[108]), .B(\round_key_gen.trw[12] ), 
         .C(\round_key_gen.trw[20] ), .D(n35834), .Z(n4_adj_8367)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)))+!A !(B (C+!(D))+!B (C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i1_4_lut_adj_544.init = 16'h5a66;
    LUT4 round_3__I_0_Mux_112_i5_3_lut (.A(\key_mem[6] [112]), .B(\key_mem[7] [112]), 
         .C(n33952), .Z(n5_adj_8368)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_112_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_87_i1_3_lut (.A(\key_mem[0] [87]), .B(\key_mem[1] [87]), 
         .C(n33952), .Z(n1_adj_8369)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_87_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_112_i4_3_lut (.A(\key_mem[4] [112]), .B(\key_mem[5] [112]), 
         .C(n33952), .Z(n4_adj_8370)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_112_i4_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_545 (.A(n33860), .B(n33640), .C(n16147), .D(n35835), 
         .Z(n16149)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_4_lut_adj_545.init = 16'ha088;
    LUT4 i10553_4_lut (.A(\key_reg[6] [13]), .B(prev_key0_reg[45]), .C(n33859), 
         .D(n33641), .Z(n16147)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i10553_4_lut.init = 16'h3aca;
    LUT4 round_3__I_0_Mux_112_i2_3_lut (.A(\key_mem[2] [112]), .B(\key_mem[3] [112]), 
         .C(n33952), .Z(n2_adj_8371)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_112_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_112_i1_3_lut (.A(\key_mem[0] [112]), .B(\key_mem[1] [112]), 
         .C(n33952), .Z(n1_adj_8372)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_112_i1_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_546 (.A(prev_key0_reg[109]), .B(\round_key_gen.trw[13] ), 
         .C(\round_key_gen.trw[21] ), .D(n35834), .Z(n4_adj_8373)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)))+!A !(B (C+!(D))+!B (C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i1_4_lut_adj_546.init = 16'h5a66;
    LUT4 round_3__I_0_Mux_111_i11_3_lut (.A(\key_mem[12] [111]), .B(\key_mem[13] [111]), 
         .C(n33952), .Z(n11_adj_8)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_111_i11_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_547 (.A(n33860), .B(n33638), .C(n16207), .D(n35835), 
         .Z(n16209)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_4_lut_adj_547.init = 16'ha088;
    LUT4 i10614_4_lut (.A(\key_reg[6] [14]), .B(prev_key0_reg[46]), .C(n33859), 
         .D(n33639), .Z(n16207)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i10614_4_lut.init = 16'h3aca;
    LUT4 round_3__I_0_Mux_111_i9_3_lut (.A(\key_mem[10] [111]), .B(\key_mem[11] [111]), 
         .C(n33952), .Z(n9_adj_8375)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_111_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_111_i8_3_lut (.A(\key_mem[8] [111]), .B(\key_mem[9] [111]), 
         .C(n33952), .Z(n8_adj_8376)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_111_i8_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_548 (.A(prev_key0_reg[110]), .B(\round_key_gen.trw[14] ), 
         .C(\round_key_gen.trw[22] ), .D(n35834), .Z(n4_adj_8377)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)))+!A !(B (C+!(D))+!B (C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i1_4_lut_adj_548.init = 16'h5a66;
    LUT4 round_3__I_0_Mux_111_i5_3_lut (.A(\key_mem[6] [111]), .B(\key_mem[7] [111]), 
         .C(n33952), .Z(n5_adj_8378)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_111_i5_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_549 (.A(n33860), .B(n33636), .C(n16267), .D(n35835), 
         .Z(n16269)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_4_lut_adj_549.init = 16'ha088;
    LUT4 round_3__I_0_Mux_111_i4_3_lut (.A(\key_mem[4] [111]), .B(\key_mem[5] [111]), 
         .C(n33952), .Z(n4_adj_8379)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_111_i4_3_lut.init = 16'hcaca;
    LUT4 i10675_4_lut (.A(\key_reg[6] [15]), .B(prev_key0_reg[47]), .C(n33859), 
         .D(n33637), .Z(n16267)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i10675_4_lut.init = 16'h3aca;
    LUT4 round_3__I_0_Mux_111_i2_3_lut (.A(\key_mem[2] [111]), .B(\key_mem[3] [111]), 
         .C(n33952), .Z(n2_adj_8380)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_111_i2_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_550 (.A(prev_key0_reg[111]), .B(\round_key_gen.trw[15] ), 
         .C(\round_key_gen.trw[23] ), .D(n35834), .Z(n4_adj_8381)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)))+!A !(B (C+!(D))+!B (C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i1_4_lut_adj_550.init = 16'h5a66;
    LUT4 round_3__I_0_Mux_111_i1_3_lut (.A(\key_mem[0] [111]), .B(\key_mem[1] [111]), 
         .C(n33952), .Z(n1_adj_8382)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_111_i1_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_551 (.A(n33860), .B(n33634), .C(n16327), .D(n35835), 
         .Z(n16329)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_4_lut_adj_551.init = 16'ha088;
    LUT4 round_3__I_0_Mux_97_i1_3_lut (.A(\key_mem[0] [97]), .B(\key_mem[1] [97]), 
         .C(n33952), .Z(n1_adj_8383)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_97_i1_3_lut.init = 16'hcaca;
    LUT4 new_sboxw_23__I_0_i25_2_lut_rep_419 (.A(\new_sboxw[16] ), .B(rcon_reg[0]), 
         .Z(n33723)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(224[13:27])
    defparam new_sboxw_23__I_0_i25_2_lut_rep_419.init = 16'h6666;
    LUT4 i2_3_lut_rep_315_4_lut (.A(\new_sboxw[16] ), .B(rcon_reg[0]), .C(prev_key1_reg[120]), 
         .D(prev_key1_reg[88]), .Z(n33619)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(224[13:27])
    defparam i2_3_lut_rep_315_4_lut.init = 16'h6996;
    LUT4 i2_4_lut_rep_652 (.A(n28850), .B(n33860), .C(\key_mem_ctrl.num_rounds[2] ), 
         .D(n33859), .Z(clk_c_enable_54)) /* synthesis lut_function=(A (B (C (D))+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam i2_4_lut_rep_652.init = 16'ha020;
    LUT4 round_3__I_0_Mux_110_i11_3_lut (.A(\key_mem[12] [110]), .B(\key_mem[13] [110]), 
         .C(n33952), .Z(n11_adj_9)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_110_i11_3_lut.init = 16'hcaca;
    LUT4 i10736_4_lut (.A(\key_reg[6] [16]), .B(prev_key0_reg[48]), .C(n33859), 
         .D(n33635), .Z(n16327)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i10736_4_lut.init = 16'h3aca;
    LUT4 round_3__I_0_Mux_110_i9_3_lut (.A(\key_mem[10] [110]), .B(\key_mem[11] [110]), 
         .C(n33952), .Z(n9_adj_8385)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_110_i9_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_552 (.A(prev_key0_reg[112]), .B(\round_key_gen.trw[16] ), 
         .C(\new_sboxw[16] ), .D(n35834), .Z(n4_adj_8386)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)))+!A !(B (C+!(D))+!B (C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i1_4_lut_adj_552.init = 16'h5a66;
    LUT4 round_3__I_0_Mux_110_i8_3_lut (.A(\key_mem[8] [110]), .B(\key_mem[9] [110]), 
         .C(n33952), .Z(n8_adj_8387)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_110_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_110_i5_3_lut (.A(\key_mem[6] [110]), .B(\key_mem[7] [110]), 
         .C(n33952), .Z(n5_adj_8388)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_110_i5_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_553 (.A(n33860), .B(n33632), .C(n16387), .D(n35835), 
         .Z(n16389)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_4_lut_adj_553.init = 16'ha088;
    LUT4 i2_3_lut_rep_420 (.A(prev_key1_reg[119]), .B(prev_key1_reg[87]), 
         .C(\round_key_gen.trw[23] ), .Z(n33724)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i2_3_lut_rep_420.init = 16'h9696;
    LUT4 i10797_4_lut (.A(\key_reg[6] [17]), .B(prev_key0_reg[49]), .C(n33859), 
         .D(n33633), .Z(n16387)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i10797_4_lut.init = 16'h3aca;
    LUT4 round_3__I_0_Mux_110_i4_3_lut (.A(\key_mem[4] [110]), .B(\key_mem[5] [110]), 
         .C(n33952), .Z(n4_adj_8389)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_110_i4_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_554 (.A(prev_key0_reg[113]), .B(\round_key_gen.trw[17] ), 
         .C(\new_sboxw[17] ), .D(n35834), .Z(n4_adj_8390)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)))+!A !(B (C+!(D))+!B (C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i1_4_lut_adj_554.init = 16'h5a66;
    LUT4 round_3__I_0_Mux_86_i11_3_lut (.A(\key_mem[12] [86]), .B(\key_mem[13] [86]), 
         .C(n33952), .Z(n11_adj_10)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_86_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_110_i2_3_lut (.A(\key_mem[2] [110]), .B(\key_mem[3] [110]), 
         .C(n33952), .Z(n2_adj_8392)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_110_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_110_i1_3_lut (.A(\key_mem[0] [110]), .B(\key_mem[1] [110]), 
         .C(n33952), .Z(n1_adj_8393)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_110_i1_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_555 (.A(n33860), .B(n33630), .C(n16447), .D(n35835), 
         .Z(n16449)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_4_lut_adj_555.init = 16'ha088;
    LUT4 i10858_4_lut (.A(\key_reg[6] [18]), .B(prev_key0_reg[50]), .C(n33859), 
         .D(n33631), .Z(n16447)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i10858_4_lut.init = 16'h3aca;
    LUT4 round_3__I_0_Mux_109_i11_3_lut (.A(\key_mem[12] [109]), .B(\key_mem[13] [109]), 
         .C(n33952), .Z(n11_adj_11)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_109_i11_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_556 (.A(prev_key0_reg[114]), .B(\round_key_gen.trw[18] ), 
         .C(\new_sboxw[18] ), .D(n35834), .Z(n4_adj_8395)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)))+!A !(B (C+!(D))+!B (C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i1_4_lut_adj_556.init = 16'h5a66;
    LUT4 round_3__I_0_Mux_109_i9_3_lut (.A(\key_mem[10] [109]), .B(\key_mem[11] [109]), 
         .C(n33952), .Z(n9_adj_8396)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_109_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_109_i8_3_lut (.A(\key_mem[8] [109]), .B(\key_mem[9] [109]), 
         .C(n33952), .Z(n8_adj_8397)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_109_i8_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_557 (.A(n33860), .B(n33628), .C(n16507), .D(n35835), 
         .Z(n16509)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_4_lut_adj_557.init = 16'ha088;
    LUT4 i5_2_lut_rep_316_4_lut (.A(prev_key1_reg[119]), .B(prev_key1_reg[87]), 
         .C(\round_key_gen.trw[23] ), .D(prev_key1_reg[55]), .Z(n33620)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i5_2_lut_rep_316_4_lut.init = 16'h6996;
    LUT4 i10919_4_lut (.A(\key_reg[6] [19]), .B(prev_key0_reg[51]), .C(n33859), 
         .D(n33629), .Z(n16507)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i10919_4_lut.init = 16'h3aca;
    LUT4 round_3__I_0_Mux_109_i5_3_lut (.A(\key_mem[6] [109]), .B(\key_mem[7] [109]), 
         .C(n33952), .Z(n5_adj_8398)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_109_i5_3_lut.init = 16'hcaca;
    LUT4 i2_4_lut_rep_653 (.A(n28850), .B(n33860), .C(\key_mem_ctrl.num_rounds[2] ), 
         .D(n33859), .Z(clk_c_enable_104)) /* synthesis lut_function=(A (B (C (D))+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam i2_4_lut_rep_653.init = 16'ha020;
    LUT4 round_3__I_0_Mux_109_i4_3_lut (.A(\key_mem[4] [109]), .B(\key_mem[5] [109]), 
         .C(n33952), .Z(n4_adj_8399)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_109_i4_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_558 (.A(prev_key0_reg[115]), .B(\round_key_gen.trw[19] ), 
         .C(\new_sboxw[19] ), .D(n35834), .Z(n4_adj_8400)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)))+!A !(B (C+!(D))+!B (C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i1_4_lut_adj_558.init = 16'h5a66;
    LUT4 round_3__I_0_Mux_109_i2_3_lut (.A(\key_mem[2] [109]), .B(\key_mem[3] [109]), 
         .C(n33952), .Z(n2_adj_8401)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_109_i2_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_559 (.A(n33860), .B(n33626), .C(n16567), .D(n35835), 
         .Z(n16569)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_4_lut_adj_559.init = 16'ha088;
    LUT4 round_3__I_0_Mux_109_i1_3_lut (.A(\key_mem[0] [109]), .B(\key_mem[1] [109]), 
         .C(n33952), .Z(n1_adj_8402)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_109_i1_3_lut.init = 16'hcaca;
    LUT4 i10980_4_lut (.A(\key_reg[6] [20]), .B(prev_key0_reg[52]), .C(n33859), 
         .D(n33627), .Z(n16567)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i10980_4_lut.init = 16'h3aca;
    LUT4 i1_4_lut_adj_560 (.A(prev_key0_reg[116]), .B(\round_key_gen.trw[20] ), 
         .C(\new_sboxw[20] ), .D(n35834), .Z(n4_adj_8403)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)))+!A !(B (C+!(D))+!B (C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i1_4_lut_adj_560.init = 16'h5a66;
    LUT4 round_3__I_0_Mux_86_i9_3_lut (.A(\key_mem[10] [86]), .B(\key_mem[11] [86]), 
         .C(n33952), .Z(n9_adj_8404)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_86_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_108_i11_3_lut (.A(\key_mem[12] [108]), .B(\key_mem[13] [108]), 
         .C(n33952), .Z(n11_adj_12)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_108_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_96_i11_3_lut (.A(\key_mem[12] [96]), .B(\key_mem[13] [96]), 
         .C(n33952), .Z(n11_adj_13)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_96_i11_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_561 (.A(n33860), .B(n33624), .C(n16627), .D(n35835), 
         .Z(n16629)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_4_lut_adj_561.init = 16'ha088;
    LUT4 round_3__I_0_Mux_108_i9_3_lut (.A(\key_mem[10] [108]), .B(\key_mem[11] [108]), 
         .C(n33952), .Z(n9_adj_8407)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_108_i9_3_lut.init = 16'hcaca;
    LUT4 i11041_4_lut (.A(\key_reg[6] [21]), .B(prev_key0_reg[53]), .C(n33859), 
         .D(n33625), .Z(n16627)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i11041_4_lut.init = 16'h3aca;
    LUT4 round_3__I_0_Mux_108_i8_3_lut (.A(\key_mem[8] [108]), .B(\key_mem[9] [108]), 
         .C(n33952), .Z(n8_adj_8408)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_108_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_86_i8_3_lut (.A(\key_mem[8] [86]), .B(\key_mem[9] [86]), 
         .C(n33952), .Z(n8_adj_8409)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_86_i8_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_562 (.A(prev_key0_reg[117]), .B(\round_key_gen.trw[21] ), 
         .C(\new_sboxw[21] ), .D(n35834), .Z(n4_adj_8410)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)))+!A !(B (C+!(D))+!B (C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i1_4_lut_adj_562.init = 16'h5a66;
    LUT4 round_3__I_0_Mux_108_i5_3_lut (.A(\key_mem[6] [108]), .B(\key_mem[7] [108]), 
         .C(n33952), .Z(n5_adj_8411)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_108_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_108_i4_3_lut (.A(\key_mem[4] [108]), .B(\key_mem[5] [108]), 
         .C(n33952), .Z(n4_adj_8412)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_108_i4_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_563 (.A(n33860), .B(n33622), .C(n16687), .D(n35835), 
         .Z(n16689)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_4_lut_adj_563.init = 16'ha088;
    LUT4 round_3__I_0_Mux_86_i5_3_lut (.A(\key_mem[6] [86]), .B(\key_mem[7] [86]), 
         .C(n33952), .Z(n5_adj_8413)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_86_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_108_i2_3_lut (.A(\key_mem[2] [108]), .B(\key_mem[3] [108]), 
         .C(n33952), .Z(n2_adj_8414)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_108_i2_3_lut.init = 16'hcaca;
    LUT4 i11102_4_lut (.A(\key_reg[6] [22]), .B(prev_key0_reg[54]), .C(n33859), 
         .D(n33623), .Z(n16687)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i11102_4_lut.init = 16'h3aca;
    LUT4 round_3__I_0_Mux_108_i1_3_lut (.A(\key_mem[0] [108]), .B(\key_mem[1] [108]), 
         .C(n33952), .Z(n1_adj_8415)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_108_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_86_i4_3_lut (.A(\key_mem[4] [86]), .B(\key_mem[5] [86]), 
         .C(n33952), .Z(n4_adj_8416)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_86_i4_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_564 (.A(prev_key0_reg[118]), .B(\round_key_gen.trw[22] ), 
         .C(\new_sboxw[22] ), .D(n35834), .Z(n4_adj_8417)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)))+!A !(B (C+!(D))+!B (C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i1_4_lut_adj_564.init = 16'h5a66;
    LUT4 round_3__I_0_Mux_107_i11_3_lut (.A(\key_mem[12] [107]), .B(\key_mem[13] [107]), 
         .C(n33952), .Z(n11_adj_14)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_107_i11_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_565 (.A(n33860), .B(n33620), .C(n16747), .D(n35835), 
         .Z(n16749)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_4_lut_adj_565.init = 16'ha088;
    LUT4 i11163_4_lut (.A(\key_reg[6] [23]), .B(prev_key0_reg[55]), .C(n33859), 
         .D(n33621), .Z(n16747)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i11163_4_lut.init = 16'h3aca;
    LUT4 round_3__I_0_Mux_107_i9_3_lut (.A(\key_mem[10] [107]), .B(\key_mem[11] [107]), 
         .C(n33952), .Z(n9_adj_8419)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_107_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_107_i8_3_lut (.A(\key_mem[8] [107]), .B(\key_mem[9] [107]), 
         .C(n33952), .Z(n8_adj_8420)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_107_i8_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_566 (.A(prev_key0_reg[119]), .B(\round_key_gen.trw[23] ), 
         .C(\new_sboxw[23] ), .D(n35834), .Z(n4_adj_8421)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)))+!A !(B (C+!(D))+!B (C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i1_4_lut_adj_566.init = 16'h5a66;
    LUT4 round_3__I_0_Mux_86_i2_3_lut (.A(\key_mem[2] [86]), .B(\key_mem[3] [86]), 
         .C(n33952), .Z(n2_adj_8422)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_86_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_107_i5_3_lut (.A(\key_mem[6] [107]), .B(\key_mem[7] [107]), 
         .C(n33952), .Z(n5_adj_8423)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_107_i5_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_567 (.A(n33860), .B(n33572), .C(n16807), .D(n35835), 
         .Z(n16809)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_4_lut_adj_567.init = 16'ha088;
    LUT4 round_3__I_0_Mux_107_i4_3_lut (.A(\key_mem[4] [107]), .B(\key_mem[5] [107]), 
         .C(n33952), .Z(n4_adj_8424)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_107_i4_3_lut.init = 16'hcaca;
    LUT4 i11224_4_lut (.A(\key_reg[6] [24]), .B(prev_key0_reg[56]), .C(n33859), 
         .D(n33573), .Z(n16807)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i11224_4_lut.init = 16'h3aca;
    LUT4 round_3__I_0_Mux_86_i1_3_lut (.A(\key_mem[0] [86]), .B(\key_mem[1] [86]), 
         .C(n33952), .Z(n1_adj_8425)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_86_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_107_i2_3_lut (.A(\key_mem[2] [107]), .B(\key_mem[3] [107]), 
         .C(n33952), .Z(n2_adj_8426)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_107_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_107_i1_3_lut (.A(\key_mem[0] [107]), .B(\key_mem[1] [107]), 
         .C(n33952), .Z(n1_adj_8427)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_107_i1_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_568 (.A(prev_key0_reg[120]), .B(n33723), .C(\round_key_gen.trw[0] ), 
         .D(n35834), .Z(n4_adj_8428)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)))+!A !(B (C+!(D))+!B (C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i1_4_lut_adj_568.init = 16'h5a66;
    LUT4 round_3__I_0_Mux_106_i11_3_lut (.A(\key_mem[12] [106]), .B(\key_mem[13] [106]), 
         .C(n33952), .Z(n11_adj_15)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_106_i11_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_569 (.A(n33860), .B(n33570), .C(n16867), .D(n35835), 
         .Z(n16869)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_4_lut_adj_569.init = 16'ha088;
    LUT4 i11285_4_lut (.A(\key_reg[6] [25]), .B(prev_key0_reg[57]), .C(n33859), 
         .D(n33571), .Z(n16867)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i11285_4_lut.init = 16'h3aca;
    LUT4 i1_4_lut_adj_570 (.A(prev_key0_reg[121]), .B(\round_key_gen.trw [25]), 
         .C(\round_key_gen.trw[1] ), .D(n35834), .Z(n4_adj_8430)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)))+!A !(B (C+!(D))+!B (C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i1_4_lut_adj_570.init = 16'h5a66;
    LUT4 round_3__I_0_Mux_85_i11_3_lut (.A(\key_mem[12] [85]), .B(\key_mem[13] [85]), 
         .C(n33952), .Z(n11_adj_16)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_85_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_106_i9_3_lut (.A(\key_mem[10] [106]), .B(\key_mem[11] [106]), 
         .C(n33952), .Z(n9_adj_8432)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_106_i9_3_lut.init = 16'hcaca;
    LUT4 i34_2_lut (.A(\rcon_logic.tmp_rcon [2]), .B(\new_sboxw[17] ), .Z(\round_key_gen.trw [25])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(110[18:27])
    defparam i34_2_lut.init = 16'h6666;
    LUT4 round_3__I_0_Mux_106_i8_3_lut (.A(\key_mem[8] [106]), .B(\key_mem[9] [106]), 
         .C(n33952), .Z(n8_adj_8433)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_106_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_106_i5_3_lut (.A(\key_mem[6] [106]), .B(\key_mem[7] [106]), 
         .C(n33952), .Z(n5_adj_8434)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_106_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_106_i4_3_lut (.A(\key_mem[4] [106]), .B(\key_mem[5] [106]), 
         .C(n33952), .Z(n4_adj_8435)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_106_i4_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_571 (.A(n33860), .B(n33569), .C(n16927), .D(n35835), 
         .Z(n16929)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_4_lut_adj_571.init = 16'ha088;
    LUT4 i11346_4_lut (.A(\key_reg[6] [26]), .B(prev_key0_reg[58]), .C(n33859), 
         .D(n33568), .Z(n16927)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i11346_4_lut.init = 16'h3aca;
    LUT4 round_3__I_0_Mux_85_i9_3_lut (.A(\key_mem[10] [85]), .B(\key_mem[11] [85]), 
         .C(n33952), .Z(n9_adj_8436)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_85_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_106_i2_3_lut (.A(\key_mem[2] [106]), .B(\key_mem[3] [106]), 
         .C(n33952), .Z(n2_adj_8437)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_106_i2_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_572 (.A(prev_key0_reg[122]), .B(n33721), .C(\round_key_gen.trw[2] ), 
         .D(n35834), .Z(n4_adj_8438)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)))+!A !(B (C+!(D))+!B (C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i1_4_lut_adj_572.init = 16'h5a66;
    LUT4 round_3__I_0_Mux_106_i1_3_lut (.A(\key_mem[0] [106]), .B(\key_mem[1] [106]), 
         .C(n33952), .Z(n1_adj_8439)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_106_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_85_i8_3_lut (.A(\key_mem[8] [85]), .B(\key_mem[9] [85]), 
         .C(n33952), .Z(n8_adj_8440)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_85_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_105_i11_3_lut (.A(\key_mem[12] [105]), .B(\key_mem[13] [105]), 
         .C(n33952), .Z(n11_adj_17)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_105_i11_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_573 (.A(n33860), .B(n33566), .C(n16987), .D(n35835), 
         .Z(n16989)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_4_lut_adj_573.init = 16'ha088;
    LUT4 i11407_4_lut (.A(\key_reg[6] [27]), .B(prev_key0_reg[59]), .C(n33859), 
         .D(n33567), .Z(n16987)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i11407_4_lut.init = 16'h3aca;
    LUT4 round_3__I_0_Mux_105_i9_3_lut (.A(\key_mem[10] [105]), .B(\key_mem[11] [105]), 
         .C(n33952), .Z(n9_adj_8442)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_105_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_105_i8_3_lut (.A(\key_mem[8] [105]), .B(\key_mem[9] [105]), 
         .C(n33952), .Z(n8_adj_8443)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_105_i8_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_574 (.A(prev_key0_reg[123]), .B(n33720), .C(\round_key_gen.trw[3] ), 
         .D(n35834), .Z(n4_adj_8444)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)))+!A !(B (C+!(D))+!B (C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i1_4_lut_adj_574.init = 16'h5a66;
    LUT4 round_3__I_0_Mux_85_i5_3_lut (.A(\key_mem[6] [85]), .B(\key_mem[7] [85]), 
         .C(n33952), .Z(n5_adj_8445)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_85_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_105_i5_3_lut (.A(\key_mem[6] [105]), .B(\key_mem[7] [105]), 
         .C(n33952), .Z(n5_adj_8446)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_105_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_85_i4_3_lut (.A(\key_mem[4] [85]), .B(\key_mem[5] [85]), 
         .C(n33952), .Z(n4_adj_8447)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_85_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_105_i4_3_lut (.A(\key_mem[4] [105]), .B(\key_mem[5] [105]), 
         .C(n33952), .Z(n4_adj_8448)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_105_i4_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_575 (.A(n33860), .B(n33564), .C(n17047), .D(n35835), 
         .Z(n17049)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_4_lut_adj_575.init = 16'ha088;
    LUT4 i11468_4_lut (.A(\key_reg[6] [28]), .B(prev_key0_reg[60]), .C(n33859), 
         .D(n33565), .Z(n17047)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i11468_4_lut.init = 16'h3aca;
    LUT4 i1_4_lut_adj_576 (.A(prev_key0_reg[124]), .B(n33719), .C(\round_key_gen.trw[4] ), 
         .D(n35834), .Z(n4_adj_8449)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)))+!A !(B (C+!(D))+!B (C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i1_4_lut_adj_576.init = 16'h5a66;
    LUT4 round_3__I_0_Mux_85_i2_3_lut (.A(\key_mem[2] [85]), .B(\key_mem[3] [85]), 
         .C(n33952), .Z(n2_adj_8450)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_85_i2_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_577 (.A(n33860), .B(n33563), .C(n17107), .D(n35835), 
         .Z(n17109)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_4_lut_adj_577.init = 16'ha088;
    LUT4 i11529_4_lut (.A(\key_reg[6] [29]), .B(prev_key0_reg[61]), .C(n33859), 
         .D(n33562), .Z(n17107)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i11529_4_lut.init = 16'h3aca;
    LUT4 i1_4_lut_adj_578 (.A(prev_key0_reg[125]), .B(n33718), .C(\round_key_gen.trw[5] ), 
         .D(n35834), .Z(n4_adj_8451)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)))+!A !(B (C+!(D))+!B (C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i1_4_lut_adj_578.init = 16'h5a66;
    LUT4 round_3__I_0_Mux_85_i1_3_lut (.A(\key_mem[0] [85]), .B(\key_mem[1] [85]), 
         .C(n33952), .Z(n1_adj_8452)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_85_i1_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_579 (.A(n33860), .B(n33560), .C(n17167), .D(n35835), 
         .Z(n17169)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_4_lut_adj_579.init = 16'ha088;
    LUT4 i11590_4_lut (.A(\key_reg[6] [30]), .B(prev_key0_reg[62]), .C(n33859), 
         .D(n33561), .Z(n17167)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i11590_4_lut.init = 16'h3aca;
    LUT4 round_3__I_0_Mux_84_i11_3_lut (.A(\key_mem[12] [84]), .B(\key_mem[13] [84]), 
         .C(n33952), .Z(n11_adj_18)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_84_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_84_i9_3_lut (.A(\key_mem[10] [84]), .B(\key_mem[11] [84]), 
         .C(n33952), .Z(n9_adj_8454)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_84_i9_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_580 (.A(prev_key0_reg[126]), .B(\round_key_gen.trw [30]), 
         .C(\round_key_gen.trw[6] ), .D(n35834), .Z(n4_adj_8455)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)))+!A !(B (C+!(D))+!B (C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i1_4_lut_adj_580.init = 16'h5a66;
    LUT4 i35_2_lut (.A(\rcon_logic.tmp_rcon [7]), .B(\new_sboxw[22] ), .Z(\round_key_gen.trw [30])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(110[18:27])
    defparam i35_2_lut.init = 16'h6666;
    LUT4 i1_4_lut_adj_581 (.A(n33860), .B(n33559), .C(n17227), .D(n35835), 
         .Z(n17229)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_4_lut_adj_581.init = 16'ha088;
    LUT4 i11651_4_lut (.A(\key_reg[6] [31]), .B(prev_key0_reg[63]), .C(n33859), 
         .D(n33558), .Z(n17227)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i11651_4_lut.init = 16'h3aca;
    LUT4 round_3__I_0_Mux_84_i8_3_lut (.A(\key_mem[8] [84]), .B(\key_mem[9] [84]), 
         .C(n33952), .Z(n8_adj_8456)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_84_i8_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_582 (.A(prev_key0_reg[127]), .B(n15124), .C(\round_key_gen.trw[7] ), 
         .D(n35834), .Z(n4_adj_8457)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)))+!A !(B (C+!(D))+!B (C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i1_4_lut_adj_582.init = 16'h5a66;
    LUT4 i33_2_lut (.A(\rcon_logic.tmp_rcon [0]), .B(\new_sboxw[23] ), .Z(n15124)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(110[18:27])
    defparam i33_2_lut.init = 16'h6666;
    LUT4 round_3__I_0_Mux_84_i5_3_lut (.A(\key_mem[6] [84]), .B(\key_mem[7] [84]), 
         .C(n33952), .Z(n5_adj_8458)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_84_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_84_i4_3_lut (.A(\key_mem[4] [84]), .B(\key_mem[5] [84]), 
         .C(n33952), .Z(n4_adj_8459)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_84_i4_3_lut.init = 16'hcaca;
    LUT4 i15099_4_lut (.A(\key_reg[1] [0]), .B(n35839), .C(n8711), .D(n33860), 
         .Z(key_mem_new[64])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15099_4_lut.init = 16'hc088;
    LUT4 i3226_3_lut (.A(n33747), .B(n33557), .C(n35835), .Z(n8711)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i3226_3_lut.init = 16'hcaca;
    LUT4 i15100_4_lut (.A(\key_reg[1] [1]), .B(n35839), .C(n8713), .D(n33860), 
         .Z(key_mem_new[65])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15100_4_lut.init = 16'hc088;
    LUT4 i3228_3_lut (.A(n33746), .B(n33556), .C(n35835), .Z(n8713)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i3228_3_lut.init = 16'hcaca;
    LUT4 i15101_4_lut (.A(\key_reg[1] [2]), .B(n35839), .C(n8715), .D(n33860), 
         .Z(key_mem_new[66])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15101_4_lut.init = 16'hc088;
    LUT4 i3230_3_lut (.A(n33745), .B(n33555), .C(n35835), .Z(n8715)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i3230_3_lut.init = 16'hcaca;
    LUT4 i15102_4_lut (.A(\key_reg[1] [3]), .B(n35839), .C(n8717), .D(n33860), 
         .Z(key_mem_new[67])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15102_4_lut.init = 16'hc088;
    LUT4 round_3__I_0_Mux_84_i2_3_lut (.A(\key_mem[2] [84]), .B(\key_mem[3] [84]), 
         .C(n33952), .Z(n2_adj_8460)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_84_i2_3_lut.init = 16'hcaca;
    LUT4 i3232_3_lut (.A(n33744), .B(n33554), .C(n35835), .Z(n8717)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i3232_3_lut.init = 16'hcaca;
    LUT4 i15103_4_lut (.A(\key_reg[1] [4]), .B(n35839), .C(n8719), .D(n33860), 
         .Z(key_mem_new[68])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15103_4_lut.init = 16'hc088;
    LUT4 i3234_3_lut (.A(n33743), .B(n33553), .C(n35835), .Z(n8719)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i3234_3_lut.init = 16'hcaca;
    LUT4 i15104_4_lut (.A(\key_reg[1] [5]), .B(n35839), .C(n8721), .D(n33860), 
         .Z(key_mem_new[69])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15104_4_lut.init = 16'hc088;
    LUT4 i3236_3_lut (.A(n33742), .B(n33552), .C(n35835), .Z(n8721)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i3236_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_96_i9_3_lut (.A(\key_mem[10] [96]), .B(\key_mem[11] [96]), 
         .C(n33952), .Z(n9_adj_8461)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_96_i9_3_lut.init = 16'hcaca;
    LUT4 i6_2_lut_3_lut_adj_583 (.A(prev_key1_reg[40]), .B(n33739), .C(keymem_sboxw[8]), 
         .Z(n15837)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;
    defparam i6_2_lut_3_lut_adj_583.init = 16'h9696;
    LUT4 i2_3_lut_rep_421 (.A(prev_key1_reg[118]), .B(prev_key1_reg[86]), 
         .C(\round_key_gen.trw[22] ), .Z(n33725)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i2_3_lut_rep_421.init = 16'h9696;
    LUT4 round_3__I_0_Mux_84_i1_3_lut (.A(\key_mem[0] [84]), .B(\key_mem[1] [84]), 
         .C(n33952), .Z(n1_adj_8462)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_84_i1_3_lut.init = 16'hcaca;
    LUT4 i15105_4_lut (.A(\key_reg[1] [6]), .B(n35839), .C(n8723), .D(n33860), 
         .Z(key_mem_new[70])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15105_4_lut.init = 16'hc088;
    LUT4 i3238_3_lut (.A(n33741), .B(n33551), .C(n35835), .Z(n8723)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i3238_3_lut.init = 16'hcaca;
    LUT4 i15106_4_lut (.A(\key_reg[1] [7]), .B(n35839), .C(n8725), .D(n33860), 
         .Z(key_mem_new[71])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15106_4_lut.init = 16'hc088;
    LUT4 i3240_3_lut (.A(n33740), .B(n33550), .C(n35835), .Z(n8725)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i3240_3_lut.init = 16'hcaca;
    LUT4 i15107_4_lut (.A(\key_reg[1] [8]), .B(n35839), .C(n8727), .D(n33860), 
         .Z(key_mem_new[72])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15107_4_lut.init = 16'hc088;
    LUT4 i3242_3_lut (.A(n33739), .B(n33549), .C(n35835), .Z(n8727)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i3242_3_lut.init = 16'hcaca;
    LUT4 i15108_4_lut (.A(\key_reg[1] [9]), .B(n35839), .C(n8729), .D(n33860), 
         .Z(key_mem_new[73])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15108_4_lut.init = 16'hc088;
    LUT4 round_3__I_0_Mux_83_i11_3_lut (.A(\key_mem[12] [83]), .B(\key_mem[13] [83]), 
         .C(n33952), .Z(n11_adj_19)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_83_i11_3_lut.init = 16'hcaca;
    LUT4 i3244_3_lut (.A(n33738), .B(n33548), .C(n35835), .Z(n8729)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i3244_3_lut.init = 16'hcaca;
    LUT4 i15109_4_lut (.A(\key_reg[1] [10]), .B(n35839), .C(n8731), .D(n33860), 
         .Z(key_mem_new[74])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15109_4_lut.init = 16'hc088;
    LUT4 round_3__I_0_Mux_83_i9_3_lut (.A(\key_mem[10] [83]), .B(\key_mem[11] [83]), 
         .C(n33952), .Z(n9_adj_8464)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_83_i9_3_lut.init = 16'hcaca;
    LUT4 i3246_3_lut (.A(n33737), .B(n33547), .C(n35835), .Z(n8731)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i3246_3_lut.init = 16'hcaca;
    LUT4 i5_2_lut_rep_318_4_lut (.A(prev_key1_reg[118]), .B(prev_key1_reg[86]), 
         .C(\round_key_gen.trw[22] ), .D(prev_key1_reg[54]), .Z(n33622)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i5_2_lut_rep_318_4_lut.init = 16'h6996;
    LUT4 i15110_4_lut (.A(\key_reg[1] [11]), .B(n35839), .C(n8733), .D(n33860), 
         .Z(key_mem_new[75])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15110_4_lut.init = 16'hc088;
    LUT4 round_3__I_0_Mux_83_i8_3_lut (.A(\key_mem[8] [83]), .B(\key_mem[9] [83]), 
         .C(n33952), .Z(n8_adj_8465)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_83_i8_3_lut.init = 16'hcaca;
    LUT4 i3248_3_lut (.A(n33736), .B(n33546), .C(n35835), .Z(n8733)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i3248_3_lut.init = 16'hcaca;
    LUT4 i15111_4_lut (.A(\key_reg[1] [12]), .B(n35839), .C(n8735), .D(n33860), 
         .Z(key_mem_new[76])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15111_4_lut.init = 16'hc088;
    LUT4 round_3__I_0_Mux_83_i5_3_lut (.A(\key_mem[6] [83]), .B(\key_mem[7] [83]), 
         .C(n33952), .Z(n5_adj_8466)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_83_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_96_i8_3_lut (.A(\key_mem[8] [96]), .B(\key_mem[9] [96]), 
         .C(n33952), .Z(n8_adj_8467)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_96_i8_3_lut.init = 16'hcaca;
    LUT4 i3250_3_lut (.A(n33735), .B(n33545), .C(n35835), .Z(n8735)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i3250_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_83_i4_3_lut (.A(\key_mem[4] [83]), .B(\key_mem[5] [83]), 
         .C(n33952), .Z(n4_adj_8468)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_83_i4_3_lut.init = 16'hcaca;
    LUT4 i15112_4_lut (.A(\key_reg[1] [13]), .B(n35839), .C(n8737), .D(n33860), 
         .Z(key_mem_new[77])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15112_4_lut.init = 16'hc088;
    LUT4 i3252_3_lut (.A(n33734), .B(n33544), .C(n35835), .Z(n8737)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i3252_3_lut.init = 16'hcaca;
    LUT4 i15113_4_lut (.A(\key_reg[1] [14]), .B(n35839), .C(n8739), .D(n33860), 
         .Z(key_mem_new[78])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15113_4_lut.init = 16'hc088;
    LUT4 round_3__I_0_Mux_83_i2_3_lut (.A(\key_mem[2] [83]), .B(\key_mem[3] [83]), 
         .C(n33952), .Z(n2_adj_8469)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_83_i2_3_lut.init = 16'hcaca;
    LUT4 i3254_3_lut (.A(n33733), .B(n33543), .C(n35835), .Z(n8739)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i3254_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_83_i1_3_lut (.A(\key_mem[0] [83]), .B(\key_mem[1] [83]), 
         .C(n33952), .Z(n1_adj_8470)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_83_i1_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_rep_422 (.A(prev_key1_reg[117]), .B(prev_key1_reg[85]), 
         .C(\round_key_gen.trw[21] ), .Z(n33726)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i2_3_lut_rep_422.init = 16'h9696;
    LUT4 round_3__I_0_Mux_96_i5_3_lut (.A(\key_mem[6] [96]), .B(\key_mem[7] [96]), 
         .C(n33952), .Z(n5_adj_8471)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_96_i5_3_lut.init = 16'hcaca;
    LUT4 i15114_4_lut (.A(\key_reg[1] [15]), .B(n35839), .C(n8741), .D(n33860), 
         .Z(key_mem_new[79])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15114_4_lut.init = 16'hc088;
    LUT4 i3256_3_lut (.A(n33732), .B(n33542), .C(n35835), .Z(n8741)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i3256_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_96_i4_3_lut (.A(\key_mem[4] [96]), .B(\key_mem[5] [96]), 
         .C(n33952), .Z(n4_adj_8472)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_96_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_96_i2_3_lut (.A(\key_mem[2] [96]), .B(\key_mem[3] [96]), 
         .C(n33952), .Z(n2_adj_8473)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_96_i2_3_lut.init = 16'hcaca;
    LUT4 i15115_4_lut (.A(\key_reg[1] [16]), .B(n35839), .C(n8743), .D(n33860), 
         .Z(key_mem_new[80])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15115_4_lut.init = 16'hc088;
    LUT4 i2_2_lut_rep_347 (.A(prev_key0_reg[72]), .B(n4_adj_8343), .Z(n33651)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i2_2_lut_rep_347.init = 16'h6666;
    LUT4 round_3__I_0_Mux_82_i11_3_lut (.A(\key_mem[12] [82]), .B(\key_mem[13] [82]), 
         .C(n33952), .Z(n11_adj_20)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_82_i11_3_lut.init = 16'hcaca;
    LUT4 i3258_3_lut (.A(n33731), .B(n33541), .C(n35835), .Z(n8743)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i3258_3_lut.init = 16'hcaca;
    LUT4 i15116_4_lut (.A(\key_reg[1] [17]), .B(n35839), .C(n8745), .D(n33860), 
         .Z(key_mem_new[81])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15116_4_lut.init = 16'hc088;
    LUT4 i3260_3_lut (.A(n33730), .B(n33540), .C(n35835), .Z(n8745)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i3260_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_82_i9_3_lut (.A(\key_mem[10] [82]), .B(\key_mem[11] [82]), 
         .C(n33952), .Z(n9_adj_8475)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_82_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_96_i1_3_lut (.A(\key_mem[0] [96]), .B(\key_mem[1] [96]), 
         .C(n33952), .Z(n1_adj_8476)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_96_i1_3_lut.init = 16'hcaca;
    LUT4 i15117_4_lut (.A(\key_reg[1] [18]), .B(n35839), .C(n8747), .D(n33860), 
         .Z(key_mem_new[82])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15117_4_lut.init = 16'hc088;
    LUT4 round_3__I_0_Mux_82_i8_3_lut (.A(\key_mem[8] [82]), .B(\key_mem[9] [82]), 
         .C(n33952), .Z(n8_adj_8477)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_82_i8_3_lut.init = 16'hcaca;
    LUT4 i3262_3_lut (.A(n33729), .B(n33539), .C(n35835), .Z(n8747)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i3262_3_lut.init = 16'hcaca;
    LUT4 i15118_4_lut (.A(\key_reg[1] [19]), .B(n35839), .C(n8749), .D(n33860), 
         .Z(key_mem_new[83])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15118_4_lut.init = 16'hc088;
    LUT4 i3264_3_lut (.A(n33728), .B(n33538), .C(n35835), .Z(n8749)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i3264_3_lut.init = 16'hcaca;
    LUT4 i5_2_lut_rep_320_4_lut (.A(prev_key1_reg[117]), .B(prev_key1_reg[85]), 
         .C(\round_key_gen.trw[21] ), .D(prev_key1_reg[53]), .Z(n33624)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i5_2_lut_rep_320_4_lut.init = 16'h6996;
    LUT4 round_3__I_0_Mux_82_i5_3_lut (.A(\key_mem[6] [82]), .B(\key_mem[7] [82]), 
         .C(n33952), .Z(n5_adj_8478)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_82_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_82_i4_3_lut (.A(\key_mem[4] [82]), .B(\key_mem[5] [82]), 
         .C(n33952), .Z(n4_adj_8479)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_82_i4_3_lut.init = 16'hcaca;
    LUT4 i15119_4_lut (.A(\key_reg[1] [20]), .B(n35839), .C(n8751), .D(n33860), 
         .Z(key_mem_new[84])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15119_4_lut.init = 16'hc088;
    LUT4 i3266_3_lut (.A(n33727), .B(n33537), .C(n35835), .Z(n8751)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i3266_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_82_i2_3_lut (.A(\key_mem[2] [82]), .B(\key_mem[3] [82]), 
         .C(n33952), .Z(n2_adj_8480)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_82_i2_3_lut.init = 16'hcaca;
    LUT4 i15120_4_lut (.A(\key_reg[1] [21]), .B(n35839), .C(n8753), .D(n33860), 
         .Z(key_mem_new[85])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15120_4_lut.init = 16'hc088;
    LUT4 i3268_3_lut (.A(n33726), .B(n33536), .C(n35835), .Z(n8753)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i3268_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_82_i1_3_lut (.A(\key_mem[0] [82]), .B(\key_mem[1] [82]), 
         .C(n33952), .Z(n1_adj_8481)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_82_i1_3_lut.init = 16'hcaca;
    LUT4 i15121_4_lut (.A(\key_reg[1] [22]), .B(n35839), .C(n8755), .D(n33860), 
         .Z(key_mem_new[86])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15121_4_lut.init = 16'hc088;
    LUT4 i3270_3_lut (.A(n33725), .B(n33535), .C(n35835), .Z(n8755)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i3270_3_lut.init = 16'hcaca;
    LUT4 i15122_4_lut (.A(\key_reg[1] [23]), .B(n35839), .C(n8757), .D(n33860), 
         .Z(key_mem_new[87])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15122_4_lut.init = 16'hc088;
    LUT4 i15066_2_lut_4_lut (.A(\key_reg[4] [31]), .B(n4_adj_8457), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[127])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15066_2_lut_4_lut.init = 16'hca00;
    LUT4 i3272_3_lut (.A(n33724), .B(n33534), .C(n35835), .Z(n8757)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i3272_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_81_i11_3_lut (.A(\key_mem[12] [81]), .B(\key_mem[13] [81]), 
         .C(n33952), .Z(n11_adj_21)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_81_i11_3_lut.init = 16'hcaca;
    LUT4 i15123_4_lut (.A(\key_reg[1] [24]), .B(n35839), .C(n8759), .D(n33860), 
         .Z(key_mem_new[88])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15123_4_lut.init = 16'hc088;
    LUT4 i3274_3_lut (.A(n33619), .B(n33517), .C(n35835), .Z(n8759)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i3274_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_81_i9_3_lut (.A(\key_mem[10] [81]), .B(\key_mem[11] [81]), 
         .C(n33952), .Z(n9_adj_8483)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_81_i9_3_lut.init = 16'hcaca;
    LUT4 i15124_4_lut (.A(\key_reg[1] [25]), .B(n35839), .C(n8761), .D(n33860), 
         .Z(key_mem_new[89])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15124_4_lut.init = 16'hc088;
    LUT4 round_3__I_0_Mux_81_i8_3_lut (.A(\key_mem[8] [81]), .B(\key_mem[9] [81]), 
         .C(n33952), .Z(n8_adj_8484)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_81_i8_3_lut.init = 16'hcaca;
    LUT4 i15125_4_lut (.A(\key_reg[1] [26]), .B(n35839), .C(n8763), .D(n33860), 
         .Z(key_mem_new[90])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15125_4_lut.init = 16'hc088;
    LUT4 i3278_3_lut (.A(n33618), .B(n33515), .C(n35835), .Z(n8763)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i3278_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_81_i5_3_lut (.A(\key_mem[6] [81]), .B(\key_mem[7] [81]), 
         .C(n33952), .Z(n5_adj_8485)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_81_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_81_i4_3_lut (.A(\key_mem[4] [81]), .B(\key_mem[5] [81]), 
         .C(n33952), .Z(n4_adj_8486)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_81_i4_3_lut.init = 16'hcaca;
    LUT4 i15126_4_lut (.A(\key_reg[1] [27]), .B(n35839), .C(n8765), .D(n33860), 
         .Z(key_mem_new[91])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15126_4_lut.init = 16'hc088;
    LUT4 i3280_3_lut (.A(n33617), .B(n33514), .C(n35835), .Z(n8765)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i3280_3_lut.init = 16'hcaca;
    LUT4 i15127_4_lut (.A(\key_reg[1] [28]), .B(n35839), .C(n8767), .D(n33860), 
         .Z(key_mem_new[92])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15127_4_lut.init = 16'hc088;
    LUT4 round_3__I_0_Mux_81_i2_3_lut (.A(\key_mem[2] [81]), .B(\key_mem[3] [81]), 
         .C(n33952), .Z(n2_adj_8487)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_81_i2_3_lut.init = 16'hcaca;
    LUT4 i3282_3_lut (.A(n33616), .B(n33513), .C(n35835), .Z(n8767)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i3282_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_81_i1_3_lut (.A(\key_mem[0] [81]), .B(\key_mem[1] [81]), 
         .C(n33952), .Z(n1_adj_8488)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_81_i1_3_lut.init = 16'hcaca;
    LUT4 i15128_4_lut (.A(\key_reg[1] [29]), .B(n35839), .C(n8769), .D(n33860), 
         .Z(key_mem_new[93])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15128_4_lut.init = 16'hc088;
    LUT4 i3284_3_lut (.A(n33615), .B(n33512), .C(n35835), .Z(n8769)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i3284_3_lut.init = 16'hcaca;
    LUT4 i15129_4_lut (.A(\key_reg[1] [30]), .B(n35839), .C(n8771), .D(n33860), 
         .Z(key_mem_new[94])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15129_4_lut.init = 16'hc088;
    LUT4 round_3__I_0_Mux_80_i11_3_lut (.A(\key_mem[12] [80]), .B(\key_mem[13] [80]), 
         .C(n33952), .Z(n11_adj_22)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_80_i11_3_lut.init = 16'hcaca;
    LUT4 i15130_4_lut (.A(\key_reg[1] [31]), .B(n35839), .C(n8773), .D(n33860), 
         .Z(key_mem_new[95])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15130_4_lut.init = 16'hc088;
    LUT4 round_3__I_0_Mux_95_i11_3_lut (.A(\key_mem[12] [95]), .B(\key_mem[13] [95]), 
         .C(n33952), .Z(n11_adj_23)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_95_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_80_i9_3_lut (.A(\key_mem[10] [80]), .B(\key_mem[11] [80]), 
         .C(n33952), .Z(n9_adj_8491)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_80_i9_3_lut.init = 16'hcaca;
    LUT4 i15131_4_lut (.A(\key_reg[0] [0]), .B(n35839), .C(n8775), .D(n33860), 
         .Z(key_mem_new[96])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15131_4_lut.init = 16'hc088;
    LUT4 round_3__I_0_Mux_80_i8_3_lut (.A(\key_mem[8] [80]), .B(\key_mem[9] [80]), 
         .C(n33952), .Z(n8_adj_8492)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_80_i8_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_rep_423 (.A(prev_key1_reg[116]), .B(prev_key1_reg[84]), 
         .C(\round_key_gen.trw[20] ), .Z(n33727)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i2_3_lut_rep_423.init = 16'h9696;
    LUT4 i15132_4_lut (.A(\key_reg[0] [1]), .B(n35839), .C(n8777), .D(n33860), 
         .Z(key_mem_new[97])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15132_4_lut.init = 16'hc088;
    LUT4 round_3__I_0_Mux_80_i5_3_lut (.A(\key_mem[6] [80]), .B(\key_mem[7] [80]), 
         .C(n33952), .Z(n5_adj_8493)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_80_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_80_i4_3_lut (.A(\key_mem[4] [80]), .B(\key_mem[5] [80]), 
         .C(n33952), .Z(n4_adj_8494)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_80_i4_3_lut.init = 16'hcaca;
    LUT4 i15133_4_lut (.A(\key_reg[0] [2]), .B(n35839), .C(n8779), .D(n33860), 
         .Z(key_mem_new[98])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15133_4_lut.init = 16'hc088;
    LUT4 round_3__I_0_Mux_80_i2_3_lut (.A(\key_mem[2] [80]), .B(\key_mem[3] [80]), 
         .C(n33952), .Z(n2_adj_8495)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_80_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_80_i1_3_lut (.A(\key_mem[0] [80]), .B(\key_mem[1] [80]), 
         .C(n33952), .Z(n1_adj_8496)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_80_i1_3_lut.init = 16'hcaca;
    LUT4 i15134_4_lut (.A(\key_reg[0] [3]), .B(n35839), .C(n8781), .D(n33860), 
         .Z(key_mem_new[99])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15134_4_lut.init = 16'hc088;
    LUT4 i15135_4_lut (.A(\key_reg[0] [4]), .B(n35839), .C(n8783), .D(n33860), 
         .Z(key_mem_new[100])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15135_4_lut.init = 16'hc088;
    LUT4 i15136_4_lut (.A(\key_reg[0] [5]), .B(n35839), .C(n8785), .D(n33860), 
         .Z(key_mem_new[101])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15136_4_lut.init = 16'hc088;
    LUT4 round_3__I_0_Mux_79_i11_3_lut (.A(\key_mem[12] [79]), .B(\key_mem[13] [79]), 
         .C(n33952), .Z(n11_adj_24)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_79_i11_3_lut.init = 16'hcaca;
    LUT4 i15137_4_lut (.A(\key_reg[0] [6]), .B(n35839), .C(n8787), .D(n33860), 
         .Z(key_mem_new[102])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15137_4_lut.init = 16'hc088;
    LUT4 i15138_4_lut (.A(\key_reg[0] [7]), .B(n35839), .C(n8789), .D(n33860), 
         .Z(key_mem_new[103])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15138_4_lut.init = 16'hc088;
    LUT4 round_3__I_0_Mux_79_i9_3_lut (.A(\key_mem[10] [79]), .B(\key_mem[11] [79]), 
         .C(n33952), .Z(n9_adj_8498)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_79_i9_3_lut.init = 16'hcaca;
    LUT4 i15139_4_lut (.A(\key_reg[0] [8]), .B(n35839), .C(n8791), .D(n33860), 
         .Z(key_mem_new[104])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15139_4_lut.init = 16'hc088;
    LUT4 round_3__I_0_Mux_79_i8_3_lut (.A(\key_mem[8] [79]), .B(\key_mem[9] [79]), 
         .C(n33952), .Z(n8_adj_8499)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_79_i8_3_lut.init = 16'hcaca;
    LUT4 i5_2_lut_rep_322_4_lut (.A(prev_key1_reg[116]), .B(prev_key1_reg[84]), 
         .C(\round_key_gen.trw[20] ), .D(prev_key1_reg[52]), .Z(n33626)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i5_2_lut_rep_322_4_lut.init = 16'h6996;
    LUT4 i15140_4_lut (.A(\key_reg[0] [9]), .B(n35839), .C(n8793), .D(n33860), 
         .Z(key_mem_new[105])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15140_4_lut.init = 16'hc088;
    LUT4 i2_3_lut_rep_424 (.A(prev_key1_reg[115]), .B(prev_key1_reg[83]), 
         .C(\round_key_gen.trw[19] ), .Z(n33728)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i2_3_lut_rep_424.init = 16'h9696;
    LUT4 round_3__I_0_Mux_79_i5_3_lut (.A(\key_mem[6] [79]), .B(\key_mem[7] [79]), 
         .C(n33952), .Z(n5_adj_8500)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_79_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_79_i4_3_lut (.A(\key_mem[4] [79]), .B(\key_mem[5] [79]), 
         .C(n33952), .Z(n4_adj_8501)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_79_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_95_i9_3_lut (.A(\key_mem[10] [95]), .B(\key_mem[11] [95]), 
         .C(n33952), .Z(n9_adj_8502)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_95_i9_3_lut.init = 16'hcaca;
    LUT4 i15141_4_lut (.A(\key_reg[0] [10]), .B(n35839), .C(n8795), .D(n33860), 
         .Z(key_mem_new[106])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15141_4_lut.init = 16'hc088;
    LUT4 i15142_4_lut (.A(\key_reg[0] [11]), .B(n35839), .C(n8797), .D(n33860), 
         .Z(key_mem_new[107])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15142_4_lut.init = 16'hc088;
    LUT4 round_3__I_0_Mux_79_i2_3_lut (.A(\key_mem[2] [79]), .B(\key_mem[3] [79]), 
         .C(n33952), .Z(n2_adj_8503)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_79_i2_3_lut.init = 16'hcaca;
    LUT4 i15143_4_lut (.A(\key_reg[0] [12]), .B(n35839), .C(n8799), .D(n33860), 
         .Z(key_mem_new[108])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15143_4_lut.init = 16'hc088;
    LUT4 round_3__I_0_Mux_79_i1_3_lut (.A(\key_mem[0] [79]), .B(\key_mem[1] [79]), 
         .C(n33952), .Z(n1_adj_8504)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_79_i1_3_lut.init = 16'hcaca;
    LUT4 i15144_4_lut (.A(\key_reg[0] [13]), .B(n35839), .C(n8801), .D(n33860), 
         .Z(key_mem_new[109])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15144_4_lut.init = 16'hc088;
    LUT4 round_3__I_0_Mux_78_i11_3_lut (.A(\key_mem[12] [78]), .B(\key_mem[13] [78]), 
         .C(n33952), .Z(n11_adj_25)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_78_i11_3_lut.init = 16'hcaca;
    LUT4 i15145_4_lut (.A(\key_reg[0] [14]), .B(n35839), .C(n8803), .D(n33860), 
         .Z(key_mem_new[110])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15145_4_lut.init = 16'hc088;
    LUT4 i15146_4_lut (.A(\key_reg[0] [15]), .B(n35839), .C(n8805), .D(n33860), 
         .Z(key_mem_new[111])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15146_4_lut.init = 16'hc088;
    LUT4 round_3__I_0_Mux_78_i9_3_lut (.A(\key_mem[10] [78]), .B(\key_mem[11] [78]), 
         .C(n33952), .Z(n9_adj_8506)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_78_i9_3_lut.init = 16'hcaca;
    LUT4 i15147_4_lut (.A(\key_reg[0] [16]), .B(n35839), .C(n8807), .D(n33860), 
         .Z(key_mem_new[112])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15147_4_lut.init = 16'hc088;
    LUT4 i15148_4_lut (.A(\key_reg[0] [17]), .B(n35839), .C(n8809), .D(n33860), 
         .Z(key_mem_new[113])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15148_4_lut.init = 16'hc088;
    LUT4 round_3__I_0_Mux_78_i8_3_lut (.A(\key_mem[8] [78]), .B(\key_mem[9] [78]), 
         .C(n33952), .Z(n8_adj_8507)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_78_i8_3_lut.init = 16'hcaca;
    LUT4 i15149_4_lut (.A(\key_reg[0] [18]), .B(n35839), .C(n8811), .D(n33860), 
         .Z(key_mem_new[114])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15149_4_lut.init = 16'hc088;
    LUT4 round_3__I_0_Mux_95_i8_3_lut (.A(\key_mem[8] [95]), .B(\key_mem[9] [95]), 
         .C(n33952), .Z(n8_adj_8508)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_95_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_78_i5_3_lut (.A(\key_mem[6] [78]), .B(\key_mem[7] [78]), 
         .C(n33952), .Z(n5_adj_8509)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_78_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_78_i4_3_lut (.A(\key_mem[4] [78]), .B(\key_mem[5] [78]), 
         .C(n33952), .Z(n4_adj_8510)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_78_i4_3_lut.init = 16'hcaca;
    LUT4 i15150_4_lut (.A(\key_reg[0] [19]), .B(n35839), .C(n8813), .D(n33860), 
         .Z(key_mem_new[115])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15150_4_lut.init = 16'hc088;
    LUT4 round_3__I_0_Mux_78_i2_3_lut (.A(\key_mem[2] [78]), .B(\key_mem[3] [78]), 
         .C(n33952), .Z(n2_adj_8511)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_78_i2_3_lut.init = 16'hcaca;
    LUT4 i15151_4_lut (.A(\key_reg[0] [20]), .B(n35839), .C(n8815), .D(n33860), 
         .Z(key_mem_new[116])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15151_4_lut.init = 16'hc088;
    LUT4 mux_85_i73_3_lut_rep_245_4_lut (.A(prev_key0_reg[72]), .B(n4_adj_8343), 
         .C(n33859), .D(\key_reg[5] [8]), .Z(n33549)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam mux_85_i73_3_lut_rep_245_4_lut.init = 16'h6f60;
    LUT4 i15152_4_lut (.A(\key_reg[0] [21]), .B(n35839), .C(n8817), .D(n33860), 
         .Z(key_mem_new[117])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15152_4_lut.init = 16'hc088;
    LUT4 round_3__I_0_Mux_78_i1_3_lut (.A(\key_mem[0] [78]), .B(\key_mem[1] [78]), 
         .C(n33952), .Z(n1_adj_8512)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_78_i1_3_lut.init = 16'hcaca;
    LUT4 i15153_4_lut (.A(\key_reg[0] [22]), .B(n35839), .C(n8819), .D(n33860), 
         .Z(key_mem_new[118])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15153_4_lut.init = 16'hc088;
    LUT4 i15154_4_lut (.A(\key_reg[0] [23]), .B(n35839), .C(n8821), .D(n33860), 
         .Z(key_mem_new[119])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15154_4_lut.init = 16'hc088;
    LUT4 round_3__I_0_Mux_77_i11_3_lut (.A(\key_mem[12] [77]), .B(\key_mem[13] [77]), 
         .C(n33952), .Z(n11_adj_26)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_77_i11_3_lut.init = 16'hcaca;
    LUT4 i15155_4_lut (.A(\key_reg[0] [24]), .B(n35839), .C(n8823), .D(n33860), 
         .Z(key_mem_new[120])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15155_4_lut.init = 16'hc088;
    LUT4 i15156_4_lut (.A(\key_reg[0] [25]), .B(n35839), .C(n8825), .D(n33860), 
         .Z(key_mem_new[121])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15156_4_lut.init = 16'hc088;
    LUT4 round_3__I_0_Mux_77_i9_3_lut (.A(\key_mem[10] [77]), .B(\key_mem[11] [77]), 
         .C(n33952), .Z(n9_adj_8514)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_77_i9_3_lut.init = 16'hcaca;
    LUT4 i3340_3_lut (.A(n33722), .B(n33532), .C(n35835), .Z(n8825)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i3340_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_77_i8_3_lut (.A(\key_mem[8] [77]), .B(\key_mem[9] [77]), 
         .C(n33952), .Z(n8_adj_8515)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_77_i8_3_lut.init = 16'hcaca;
    LUT4 i15157_4_lut (.A(\key_reg[0] [26]), .B(n35839), .C(n8827), .D(n33860), 
         .Z(key_mem_new[122])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15157_4_lut.init = 16'hc088;
    LUT4 i15158_4_lut (.A(\key_reg[0] [27]), .B(n35839), .C(n8829), .D(n33860), 
         .Z(key_mem_new[123])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15158_4_lut.init = 16'hc088;
    LUT4 i15159_4_lut (.A(\key_reg[0] [28]), .B(n35839), .C(n8831), .D(n33860), 
         .Z(key_mem_new[124])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15159_4_lut.init = 16'hc088;
    LUT4 round_3__I_0_Mux_77_i5_3_lut (.A(\key_mem[6] [77]), .B(\key_mem[7] [77]), 
         .C(n33952), .Z(n5_adj_8516)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_77_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_77_i4_3_lut (.A(\key_mem[4] [77]), .B(\key_mem[5] [77]), 
         .C(n33952), .Z(n4_adj_8517)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_77_i4_3_lut.init = 16'hcaca;
    LUT4 i15160_4_lut (.A(\key_reg[0] [29]), .B(n35839), .C(n8833), .D(n33860), 
         .Z(key_mem_new[125])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15160_4_lut.init = 16'hc088;
    LUT4 round_3__I_0_Mux_77_i2_3_lut (.A(\key_mem[2] [77]), .B(\key_mem[3] [77]), 
         .C(n33952), .Z(n2_adj_8518)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_77_i2_3_lut.init = 16'hcaca;
    LUT4 i15161_4_lut (.A(\key_reg[0] [30]), .B(n35839), .C(n8835), .D(n33860), 
         .Z(key_mem_new[126])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15161_4_lut.init = 16'hc088;
    LUT4 i3350_3_lut (.A(n33717), .B(n33527), .C(n35835), .Z(n8835)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i3350_3_lut.init = 16'hcaca;
    LUT4 i15162_4_lut (.A(\key_reg[0] [31]), .B(n35839), .C(n8837), .D(n33860), 
         .Z(key_mem_new[127])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(228[7] 302[12])
    defparam i15162_4_lut.init = 16'hc088;
    LUT4 i3352_3_lut (.A(n33716), .B(n33526), .C(n35835), .Z(n8837)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(232[11] 301[18])
    defparam i3352_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_77_i1_3_lut (.A(\key_mem[0] [77]), .B(\key_mem[1] [77]), 
         .C(n33952), .Z(n1_adj_8519)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_77_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_76_i11_3_lut (.A(\key_mem[12] [76]), .B(\key_mem[13] [76]), 
         .C(n33952), .Z(n11_adj_27)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_76_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_76_i9_3_lut (.A(\key_mem[10] [76]), .B(\key_mem[11] [76]), 
         .C(n33952), .Z(n9_adj_8521)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_76_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_76_i8_3_lut (.A(\key_mem[8] [76]), .B(\key_mem[9] [76]), 
         .C(n33952), .Z(n8_adj_8522)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_76_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_76_i5_3_lut (.A(\key_mem[6] [76]), .B(\key_mem[7] [76]), 
         .C(n33952), .Z(n5_adj_8523)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_76_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_76_i4_3_lut (.A(\key_mem[4] [76]), .B(\key_mem[5] [76]), 
         .C(n33952), .Z(n4_adj_8524)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_76_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_76_i2_3_lut (.A(\key_mem[2] [76]), .B(\key_mem[3] [76]), 
         .C(n33952), .Z(n2_adj_8525)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_76_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_76_i1_3_lut (.A(\key_mem[0] [76]), .B(\key_mem[1] [76]), 
         .C(n33952), .Z(n1_adj_8526)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_76_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_75_i11_3_lut (.A(\key_mem[12] [75]), .B(\key_mem[13] [75]), 
         .C(n33952), .Z(n11_adj_28)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_75_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_75_i9_3_lut (.A(\key_mem[10] [75]), .B(\key_mem[11] [75]), 
         .C(n33952), .Z(n9_adj_8528)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_75_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_75_i8_3_lut (.A(\key_mem[8] [75]), .B(\key_mem[9] [75]), 
         .C(n33952), .Z(n8_adj_8529)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_75_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_75_i5_3_lut (.A(\key_mem[6] [75]), .B(\key_mem[7] [75]), 
         .C(n33952), .Z(n5_adj_8530)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_75_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_75_i4_3_lut (.A(\key_mem[4] [75]), .B(\key_mem[5] [75]), 
         .C(n33952), .Z(n4_adj_8531)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_75_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_75_i2_3_lut (.A(\key_mem[2] [75]), .B(\key_mem[3] [75]), 
         .C(n33952), .Z(n2_adj_8532)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_75_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_75_i1_3_lut (.A(\key_mem[0] [75]), .B(\key_mem[1] [75]), 
         .C(n33952), .Z(n1_adj_8533)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_75_i1_3_lut.init = 16'hcaca;
    LUT4 i5_2_lut_rep_324_4_lut (.A(prev_key1_reg[115]), .B(prev_key1_reg[83]), 
         .C(\round_key_gen.trw[19] ), .D(prev_key1_reg[51]), .Z(n33628)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i5_2_lut_rep_324_4_lut.init = 16'h6996;
    LUT4 i2_3_lut_rep_425 (.A(prev_key1_reg[114]), .B(prev_key1_reg[82]), 
         .C(\round_key_gen.trw[18] ), .Z(n33729)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i2_3_lut_rep_425.init = 16'h9696;
    LUT4 round_3__I_0_Mux_74_i11_3_lut (.A(\key_mem[12] [74]), .B(\key_mem[13] [74]), 
         .C(n33952), .Z(n11_adj_29)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_74_i11_3_lut.init = 16'hcaca;
    LUT4 i15065_2_lut_4_lut (.A(\key_reg[4] [30]), .B(n4_adj_8455), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[126])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15065_2_lut_4_lut.init = 16'hca00;
    LUT4 round_3__I_0_Mux_95_i5_3_lut (.A(\key_mem[6] [95]), .B(\key_mem[7] [95]), 
         .C(n33952), .Z(n5_adj_8535)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_95_i5_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut (.A(n35839), .B(n72), .Z(rcon_we)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam i1_2_lut.init = 16'hdddd;
    LUT4 round_3__I_0_Mux_95_i4_3_lut (.A(\key_mem[4] [95]), .B(\key_mem[5] [95]), 
         .C(n33952), .Z(n4_adj_8536)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_95_i4_3_lut.init = 16'hcaca;
    LUT4 i15033_2_lut_4_lut (.A(\key_reg[5] [30]), .B(n33561), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[94])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15033_2_lut_4_lut.init = 16'hca00;
    LUT4 round_3__I_0_Mux_74_i9_3_lut (.A(\key_mem[10] [74]), .B(\key_mem[11] [74]), 
         .C(n33952), .Z(n9_adj_8537)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_74_i9_3_lut.init = 16'hcaca;
    LUT4 i5_2_lut_rep_326_4_lut (.A(prev_key1_reg[114]), .B(prev_key1_reg[82]), 
         .C(\round_key_gen.trw[18] ), .D(prev_key1_reg[50]), .Z(n33630)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i5_2_lut_rep_326_4_lut.init = 16'h6996;
    LUT4 round_3__I_0_Mux_74_i8_3_lut (.A(\key_mem[8] [74]), .B(\key_mem[9] [74]), 
         .C(n33952), .Z(n8_adj_8538)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_74_i8_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_adj_584 (.A(n35839), .B(\rcon_logic.tmp_rcon [0]), .C(n72), 
         .Z(rcon_new[0])) /* synthesis lut_function=((B (C))+!A) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam i1_3_lut_adj_584.init = 16'hd5d5;
    LUT4 round_3__I_0_Mux_74_i5_3_lut (.A(\key_mem[6] [74]), .B(\key_mem[7] [74]), 
         .C(n33952), .Z(n5_adj_8539)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_74_i5_3_lut.init = 16'hcaca;
    LUT4 i15032_2_lut_4_lut (.A(\key_reg[5] [29]), .B(n33562), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[93])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15032_2_lut_4_lut.init = 16'hca00;
    LUT4 round_3__I_0_Mux_74_i4_3_lut (.A(\key_mem[4] [74]), .B(\key_mem[5] [74]), 
         .C(n33952), .Z(n4_adj_8540)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_74_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_74_i2_3_lut (.A(\key_mem[2] [74]), .B(\key_mem[3] [74]), 
         .C(n33952), .Z(n2_adj_8541)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_74_i2_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_rep_426 (.A(prev_key1_reg[113]), .B(prev_key1_reg[81]), 
         .C(\round_key_gen.trw[17] ), .Z(n33730)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i2_3_lut_rep_426.init = 16'h9696;
    LUT4 i1_4_lut_adj_585 (.A(n33860), .B(\key_mem_ctrl.num_rounds[2] ), 
         .C(n33859), .D(n35834), .Z(n72)) /* synthesis lut_function=(A (((D)+!C)+!B)+!A !(B)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam i1_4_lut_adj_585.init = 16'hbb3b;
    LUT4 i6_2_lut_3_lut_adj_586 (.A(prev_key1_reg[39]), .B(n33740), .C(keymem_sboxw[7]), 
         .Z(n15777)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;
    defparam i6_2_lut_3_lut_adj_586.init = 16'h9696;
    LUT4 round_3__I_0_Mux_95_i2_3_lut (.A(\key_mem[2] [95]), .B(\key_mem[3] [95]), 
         .C(n33952), .Z(n2_adj_8542)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_95_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_74_i1_3_lut (.A(\key_mem[0] [74]), .B(\key_mem[1] [74]), 
         .C(n33952), .Z(n1_adj_8543)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_74_i1_3_lut.init = 16'hcaca;
    LUT4 i5_2_lut_rep_328_4_lut (.A(prev_key1_reg[113]), .B(prev_key1_reg[81]), 
         .C(\round_key_gen.trw[17] ), .D(prev_key1_reg[49]), .Z(n33632)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i5_2_lut_rep_328_4_lut.init = 16'h6996;
    LUT4 i2_2_lut_rep_349 (.A(prev_key0_reg[71]), .B(n4_adj_8339), .Z(n33653)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i2_2_lut_rep_349.init = 16'h6666;
    LUT4 i15031_2_lut_4_lut (.A(\key_reg[5] [28]), .B(n33565), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[92])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15031_2_lut_4_lut.init = 16'hca00;
    LUT4 i2_3_lut_rep_427 (.A(prev_key1_reg[112]), .B(prev_key1_reg[80]), 
         .C(\round_key_gen.trw[16] ), .Z(n33731)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i2_3_lut_rep_427.init = 16'h9696;
    LUT4 round_3__I_0_Mux_73_i11_3_lut (.A(\key_mem[12] [73]), .B(\key_mem[13] [73]), 
         .C(n33952), .Z(n11_adj_30)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_73_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_95_i1_3_lut (.A(\key_mem[0] [95]), .B(\key_mem[1] [95]), 
         .C(n33952), .Z(n1_adj_8545)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_95_i1_3_lut.init = 16'hcaca;
    LUT4 i5_2_lut_rep_330_4_lut (.A(prev_key1_reg[112]), .B(prev_key1_reg[80]), 
         .C(\round_key_gen.trw[16] ), .D(prev_key1_reg[48]), .Z(n33634)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i5_2_lut_rep_330_4_lut.init = 16'h6996;
    LUT4 i15030_2_lut_4_lut (.A(\key_reg[5] [27]), .B(n33567), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[91])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15030_2_lut_4_lut.init = 16'hca00;
    LUT4 round_3__I_0_Mux_73_i9_3_lut (.A(\key_mem[10] [73]), .B(\key_mem[11] [73]), 
         .C(n33952), .Z(n9_adj_8546)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_73_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_73_i8_3_lut (.A(\key_mem[8] [73]), .B(\key_mem[9] [73]), 
         .C(n33952), .Z(n8_adj_8547)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_73_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_94_i11_3_lut (.A(\key_mem[12] [94]), .B(\key_mem[13] [94]), 
         .C(n33952), .Z(n11_adj_31)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_94_i11_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_rep_428 (.A(prev_key1_reg[111]), .B(prev_key1_reg[79]), 
         .C(\round_key_gen.trw[15] ), .Z(n33732)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i2_3_lut_rep_428.init = 16'h9696;
    LUT4 i15064_2_lut_4_lut (.A(\key_reg[4] [29]), .B(n4_adj_8451), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[125])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15064_2_lut_4_lut.init = 16'hca00;
    LUT4 round_3__I_0_Mux_94_i9_3_lut (.A(\key_mem[10] [94]), .B(\key_mem[11] [94]), 
         .C(n33952), .Z(n9_adj_8549)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_94_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_94_i8_3_lut (.A(\key_mem[8] [94]), .B(\key_mem[9] [94]), 
         .C(n33952), .Z(n8_adj_8550)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_94_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_73_i5_3_lut (.A(\key_mem[6] [73]), .B(\key_mem[7] [73]), 
         .C(n33952), .Z(n5_adj_8551)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_73_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_73_i4_3_lut (.A(\key_mem[4] [73]), .B(\key_mem[5] [73]), 
         .C(n33952), .Z(n4_adj_8552)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_73_i4_3_lut.init = 16'hcaca;
    LUT4 i5_2_lut_rep_332_4_lut (.A(prev_key1_reg[111]), .B(prev_key1_reg[79]), 
         .C(\round_key_gen.trw[15] ), .D(prev_key1_reg[47]), .Z(n33636)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i5_2_lut_rep_332_4_lut.init = 16'h6996;
    LUT4 i2_3_lut_rep_429 (.A(prev_key1_reg[110]), .B(prev_key1_reg[78]), 
         .C(\round_key_gen.trw[14] ), .Z(n33733)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i2_3_lut_rep_429.init = 16'h9696;
    LUT4 round_3__I_0_Mux_73_i2_3_lut (.A(\key_mem[2] [73]), .B(\key_mem[3] [73]), 
         .C(n33952), .Z(n2_adj_8553)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_73_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_73_i1_3_lut (.A(\key_mem[0] [73]), .B(\key_mem[1] [73]), 
         .C(n33952), .Z(n1_adj_8554)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_73_i1_3_lut.init = 16'hcaca;
    LUT4 i15029_2_lut_4_lut (.A(\key_reg[5] [26]), .B(n33568), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[90])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15029_2_lut_4_lut.init = 16'hca00;
    LUT4 round_3__I_0_Mux_94_i5_3_lut (.A(\key_mem[6] [94]), .B(\key_mem[7] [94]), 
         .C(n33952), .Z(n5_adj_8555)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_94_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_72_i11_3_lut (.A(\key_mem[12] [72]), .B(\key_mem[13] [72]), 
         .C(n33952), .Z(n11_adj_32)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_72_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_72_i9_3_lut (.A(\key_mem[10] [72]), .B(\key_mem[11] [72]), 
         .C(n33952), .Z(n9_adj_8557)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_72_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_72_i8_3_lut (.A(\key_mem[8] [72]), .B(\key_mem[9] [72]), 
         .C(n33952), .Z(n8_adj_8558)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_72_i8_3_lut.init = 16'hcaca;
    LUT4 i5_2_lut_rep_334_4_lut (.A(prev_key1_reg[110]), .B(prev_key1_reg[78]), 
         .C(\round_key_gen.trw[14] ), .D(prev_key1_reg[46]), .Z(n33638)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i5_2_lut_rep_334_4_lut.init = 16'h6996;
    LUT4 round_3__I_0_Mux_72_i5_3_lut (.A(\key_mem[6] [72]), .B(\key_mem[7] [72]), 
         .C(n33952), .Z(n5_adj_8559)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_72_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_94_i4_3_lut (.A(\key_mem[4] [94]), .B(\key_mem[5] [94]), 
         .C(n33952), .Z(n4_adj_8560)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_94_i4_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_rep_430 (.A(prev_key1_reg[109]), .B(prev_key1_reg[77]), 
         .C(\round_key_gen.trw[13] ), .Z(n33734)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i2_3_lut_rep_430.init = 16'h9696;
    LUT4 round_3__I_0_Mux_72_i4_3_lut (.A(\key_mem[4] [72]), .B(\key_mem[5] [72]), 
         .C(n33952), .Z(n4_adj_8561)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_72_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_94_i2_3_lut (.A(\key_mem[2] [94]), .B(\key_mem[3] [94]), 
         .C(n33952), .Z(n2_adj_8562)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_94_i2_3_lut.init = 16'hcaca;
    LUT4 i5_2_lut_rep_336_4_lut (.A(prev_key1_reg[109]), .B(prev_key1_reg[77]), 
         .C(\round_key_gen.trw[13] ), .D(prev_key1_reg[45]), .Z(n33640)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i5_2_lut_rep_336_4_lut.init = 16'h6996;
    LUT4 i2_3_lut_rep_431 (.A(prev_key1_reg[108]), .B(prev_key1_reg[76]), 
         .C(\round_key_gen.trw[12] ), .Z(n33735)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i2_3_lut_rep_431.init = 16'h9696;
    LUT4 round_3__I_0_Mux_94_i1_3_lut (.A(\key_mem[0] [94]), .B(\key_mem[1] [94]), 
         .C(n33952), .Z(n1_adj_8563)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_94_i1_3_lut.init = 16'hcaca;
    LUT4 i15063_2_lut_4_lut (.A(\key_reg[4] [28]), .B(n4_adj_8449), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[124])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15063_2_lut_4_lut.init = 16'hca00;
    LUT4 mux_85_i72_3_lut_rep_246_4_lut (.A(prev_key0_reg[71]), .B(n4_adj_8339), 
         .C(n33859), .D(\key_reg[5] [7]), .Z(n33550)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam mux_85_i72_3_lut_rep_246_4_lut.init = 16'h6f60;
    LUT4 i5_2_lut_rep_338_4_lut (.A(prev_key1_reg[108]), .B(prev_key1_reg[76]), 
         .C(\round_key_gen.trw[12] ), .D(prev_key1_reg[44]), .Z(n33642)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i5_2_lut_rep_338_4_lut.init = 16'h6996;
    LUT4 i2_3_lut_rep_432 (.A(prev_key1_reg[107]), .B(prev_key1_reg[75]), 
         .C(\round_key_gen.trw[11] ), .Z(n33736)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i2_3_lut_rep_432.init = 16'h9696;
    LUT4 i5_2_lut_rep_340_4_lut (.A(prev_key1_reg[107]), .B(prev_key1_reg[75]), 
         .C(\round_key_gen.trw[11] ), .D(prev_key1_reg[43]), .Z(n33644)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i5_2_lut_rep_340_4_lut.init = 16'h6996;
    LUT4 round_3__I_0_Mux_93_i11_3_lut (.A(\key_mem[12] [93]), .B(\key_mem[13] [93]), 
         .C(n33952), .Z(n11_adj_33)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_93_i11_3_lut.init = 16'hcaca;
    FD1P3AX key_mem_14___i1 (.D(key_mem_0__127__N_6752[0]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1.GSR = "ENABLED";
    FD1P3IX prev_key1_reg__i1 (.D(prev_key1_new_127__N_4787[0]), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(keymem_sboxw[0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i1.GSR = "DISABLED";
    LUT4 round_3__I_0_Mux_72_i2_3_lut (.A(\key_mem[2] [72]), .B(\key_mem[3] [72]), 
         .C(n33952), .Z(n2_adj_8565)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_72_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_72_i1_3_lut (.A(\key_mem[0] [72]), .B(\key_mem[1] [72]), 
         .C(n33952), .Z(n1_adj_8566)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_72_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_93_i9_3_lut (.A(\key_mem[10] [93]), .B(\key_mem[11] [93]), 
         .C(n33952), .Z(n9_adj_8567)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_93_i9_3_lut.init = 16'hcaca;
    LUT4 i15028_2_lut_4_lut (.A(\key_reg[5] [25]), .B(n33571), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[89])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15028_2_lut_4_lut.init = 16'hca00;
    LUT4 round_3__I_0_Mux_93_i8_3_lut (.A(\key_mem[8] [93]), .B(\key_mem[9] [93]), 
         .C(n33952), .Z(n8_adj_8568)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_93_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_71_i11_3_lut (.A(\key_mem[12] [71]), .B(\key_mem[13] [71]), 
         .C(n33952), .Z(n11_adj_34)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_71_i11_3_lut.init = 16'hcaca;
    LUT4 i11_4_lut (.A(n5), .B(keymem_sboxw[0]), .C(init_state), .D(n10), 
         .Z(muxed_sboxw[0])) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(181[17:28])
    defparam i11_4_lut.init = 16'hc5c0;
    LUT4 round_3__I_0_Mux_71_i9_3_lut (.A(\key_mem[10] [71]), .B(\key_mem[11] [71]), 
         .C(n33952), .Z(n9_adj_8571)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_71_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_71_i8_3_lut (.A(\key_mem[8] [71]), .B(\key_mem[9] [71]), 
         .C(n33952), .Z(n8_adj_8572)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_71_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_71_i5_3_lut (.A(\key_mem[6] [71]), .B(\key_mem[7] [71]), 
         .C(n33952), .Z(n5_adj_8573)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_71_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_71_i4_3_lut (.A(\key_mem[4] [71]), .B(\key_mem[5] [71]), 
         .C(n33952), .Z(n4_adj_8574)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_71_i4_3_lut.init = 16'hcaca;
    LUT4 i6_2_lut_3_lut_adj_587 (.A(prev_key1_reg[38]), .B(n33741), .C(keymem_sboxw[6]), 
         .Z(n15717)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;
    defparam i6_2_lut_3_lut_adj_587.init = 16'h9696;
    LUT4 i15027_2_lut_4_lut (.A(\key_reg[5] [24]), .B(n33573), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[88])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15027_2_lut_4_lut.init = 16'hca00;
    LUT4 round_3__I_0_Mux_71_i2_3_lut (.A(\key_mem[2] [71]), .B(\key_mem[3] [71]), 
         .C(n33952), .Z(n2_adj_8575)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_71_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_71_i1_3_lut (.A(\key_mem[0] [71]), .B(\key_mem[1] [71]), 
         .C(n33952), .Z(n1_adj_8576)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_71_i1_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_rep_433 (.A(prev_key1_reg[106]), .B(prev_key1_reg[74]), 
         .C(\round_key_gen.trw[10] ), .Z(n33737)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i2_3_lut_rep_433.init = 16'h9696;
    LUT4 i15021_2_lut_4_lut (.A(\key_reg[5] [18]), .B(n33631), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[82])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15021_2_lut_4_lut.init = 16'hca00;
    LUT4 round_3__I_0_Mux_93_i5_3_lut (.A(\key_mem[6] [93]), .B(\key_mem[7] [93]), 
         .C(n33952), .Z(n5_adj_8577)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_93_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_70_i11_3_lut (.A(\key_mem[12] [70]), .B(\key_mem[13] [70]), 
         .C(n33952), .Z(n11_adj_35)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_70_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_70_i9_3_lut (.A(\key_mem[10] [70]), .B(\key_mem[11] [70]), 
         .C(n33952), .Z(n9_adj_8579)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_70_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_70_i8_3_lut (.A(\key_mem[8] [70]), .B(\key_mem[9] [70]), 
         .C(n33952), .Z(n8_adj_8580)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_70_i8_3_lut.init = 16'hcaca;
    LUT4 i5_2_lut_rep_342_4_lut (.A(prev_key1_reg[106]), .B(prev_key1_reg[74]), 
         .C(\round_key_gen.trw[10] ), .D(prev_key1_reg[42]), .Z(n33646)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i5_2_lut_rep_342_4_lut.init = 16'h6996;
    LUT4 round_3__I_0_Mux_93_i4_3_lut (.A(\key_mem[4] [93]), .B(\key_mem[5] [93]), 
         .C(n33952), .Z(n4_adj_8581)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_93_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_70_i5_3_lut (.A(\key_mem[6] [70]), .B(\key_mem[7] [70]), 
         .C(n33952), .Z(n5_adj_8582)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_70_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_70_i4_3_lut (.A(\key_mem[4] [70]), .B(\key_mem[5] [70]), 
         .C(n33952), .Z(n4_adj_8583)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_70_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_70_i2_3_lut (.A(\key_mem[2] [70]), .B(\key_mem[3] [70]), 
         .C(n33952), .Z(n2_adj_8584)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_70_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_70_i1_3_lut (.A(\key_mem[0] [70]), .B(\key_mem[1] [70]), 
         .C(n33952), .Z(n1_adj_8585)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_70_i1_3_lut.init = 16'hcaca;
    LUT4 i2_2_lut_rep_351 (.A(prev_key0_reg[70]), .B(n4_adj_8337), .Z(n33655)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i2_2_lut_rep_351.init = 16'h6666;
    LUT4 round_3__I_0_Mux_69_i11_3_lut (.A(\key_mem[12] [69]), .B(\key_mem[13] [69]), 
         .C(n33952), .Z(n11_adj_36)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_69_i11_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_rep_434 (.A(prev_key1_reg[105]), .B(prev_key1_reg[73]), 
         .C(\round_key_gen.trw[9] ), .Z(n33738)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i2_3_lut_rep_434.init = 16'h9696;
    LUT4 i11_4_lut_adj_588 (.A(n5), .B(keymem_sboxw[1]), .C(init_state), 
         .D(n10_adj_8587), .Z(muxed_sboxw[1])) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(181[17:28])
    defparam i11_4_lut_adj_588.init = 16'hc5c0;
    LUT4 i5_2_lut_rep_344_4_lut (.A(prev_key1_reg[105]), .B(prev_key1_reg[73]), 
         .C(\round_key_gen.trw[9] ), .D(prev_key1_reg[41]), .Z(n33648)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i5_2_lut_rep_344_4_lut.init = 16'h6996;
    LUT4 i2_3_lut_rep_435 (.A(prev_key1_reg[104]), .B(prev_key1_reg[72]), 
         .C(\round_key_gen.trw[8] ), .Z(n33739)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i2_3_lut_rep_435.init = 16'h9696;
    LUT4 mux_85_i71_3_lut_rep_247_4_lut (.A(prev_key0_reg[70]), .B(n4_adj_8337), 
         .C(n33859), .D(\key_reg[5] [6]), .Z(n33551)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam mux_85_i71_3_lut_rep_247_4_lut.init = 16'h6f60;
    LUT4 round_3__I_0_Mux_93_i2_3_lut (.A(\key_mem[2] [93]), .B(\key_mem[3] [93]), 
         .C(n33952), .Z(n2_adj_8588)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_93_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_93_i1_3_lut (.A(\key_mem[0] [93]), .B(\key_mem[1] [93]), 
         .C(n33952), .Z(n1_adj_8589)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_93_i1_3_lut.init = 16'hcaca;
    LUT4 i5_2_lut_rep_346_4_lut (.A(prev_key1_reg[104]), .B(prev_key1_reg[72]), 
         .C(\round_key_gen.trw[8] ), .D(prev_key1_reg[40]), .Z(n33650)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i5_2_lut_rep_346_4_lut.init = 16'h6996;
    LUT4 i11_4_lut_adj_589 (.A(n5), .B(keymem_sboxw[2]), .C(init_state), 
         .D(n10_adj_8590), .Z(muxed_sboxw[2])) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(181[17:28])
    defparam i11_4_lut_adj_589.init = 16'hc5c0;
    LUT4 round_3__I_0_Mux_69_i9_3_lut (.A(\key_mem[10] [69]), .B(\key_mem[11] [69]), 
         .C(n33952), .Z(n9_adj_8591)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_69_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_69_i8_3_lut (.A(\key_mem[8] [69]), .B(\key_mem[9] [69]), 
         .C(n33952), .Z(n8_adj_8592)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_69_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_69_i5_3_lut (.A(\key_mem[6] [69]), .B(\key_mem[7] [69]), 
         .C(n33952), .Z(n5_adj_8593)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_69_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_69_i4_3_lut (.A(\key_mem[4] [69]), .B(\key_mem[5] [69]), 
         .C(n33952), .Z(n4_adj_8594)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_69_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_69_i2_3_lut (.A(\key_mem[2] [69]), .B(\key_mem[3] [69]), 
         .C(n33952), .Z(n2_adj_8595)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_69_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_92_i11_3_lut (.A(\key_mem[12] [92]), .B(\key_mem[13] [92]), 
         .C(n33952), .Z(n11_adj_37)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_92_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_69_i1_3_lut (.A(\key_mem[0] [69]), .B(\key_mem[1] [69]), 
         .C(n33952), .Z(n1_adj_8597)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_69_i1_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_rep_436 (.A(prev_key1_reg[103]), .B(prev_key1_reg[71]), 
         .C(\round_key_gen.trw[7] ), .Z(n33740)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i2_3_lut_rep_436.init = 16'h9696;
    LUT4 i11_4_lut_adj_590 (.A(n5), .B(keymem_sboxw[3]), .C(init_state), 
         .D(n10_adj_8598), .Z(muxed_sboxw[3])) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(181[17:28])
    defparam i11_4_lut_adj_590.init = 16'hc5c0;
    LUT4 round_3__I_0_Mux_92_i9_3_lut (.A(\key_mem[10] [92]), .B(\key_mem[11] [92]), 
         .C(n33952), .Z(n9_adj_8599)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_92_i9_3_lut.init = 16'hcaca;
    LUT4 i15020_2_lut_4_lut (.A(\key_reg[5] [17]), .B(n33633), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[81])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15020_2_lut_4_lut.init = 16'hca00;
    LUT4 round_3__I_0_Mux_68_i11_3_lut (.A(\key_mem[12] [68]), .B(\key_mem[13] [68]), 
         .C(n33952), .Z(n11_adj_38)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_68_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_92_i8_3_lut (.A(\key_mem[8] [92]), .B(\key_mem[9] [92]), 
         .C(n33952), .Z(n8_adj_8601)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_92_i8_3_lut.init = 16'hcaca;
    LUT4 i5_2_lut_rep_348_4_lut (.A(prev_key1_reg[103]), .B(prev_key1_reg[71]), 
         .C(\round_key_gen.trw[7] ), .D(prev_key1_reg[39]), .Z(n33652)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i5_2_lut_rep_348_4_lut.init = 16'h6996;
    LUT4 i2_3_lut_rep_437 (.A(prev_key1_reg[102]), .B(prev_key1_reg[70]), 
         .C(\round_key_gen.trw[6] ), .Z(n33741)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i2_3_lut_rep_437.init = 16'h9696;
    LUT4 i11_4_lut_adj_591 (.A(n5), .B(keymem_sboxw[4]), .C(init_state), 
         .D(n10_adj_8602), .Z(muxed_sboxw[4])) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(181[17:28])
    defparam i11_4_lut_adj_591.init = 16'hc5c0;
    LUT4 round_3__I_0_Mux_92_i5_3_lut (.A(\key_mem[6] [92]), .B(\key_mem[7] [92]), 
         .C(n33952), .Z(n5_adj_8603)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_92_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_92_i4_3_lut (.A(\key_mem[4] [92]), .B(\key_mem[5] [92]), 
         .C(n33952), .Z(n4_adj_8604)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_92_i4_3_lut.init = 16'hcaca;
    LUT4 i6_2_lut_3_lut_adj_592 (.A(prev_key1_reg[37]), .B(n33742), .C(keymem_sboxw[5]), 
         .Z(n15657)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;
    defparam i6_2_lut_3_lut_adj_592.init = 16'h9696;
    LUT4 round_3__I_0_Mux_68_i9_3_lut (.A(\key_mem[10] [68]), .B(\key_mem[11] [68]), 
         .C(n33952), .Z(n9_adj_8605)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_68_i9_3_lut.init = 16'hcaca;
    LUT4 i5_2_lut_rep_350_4_lut (.A(prev_key1_reg[102]), .B(prev_key1_reg[70]), 
         .C(\round_key_gen.trw[6] ), .D(prev_key1_reg[38]), .Z(n33654)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i5_2_lut_rep_350_4_lut.init = 16'h6996;
    LUT4 round_3__I_0_Mux_68_i8_3_lut (.A(\key_mem[8] [68]), .B(\key_mem[9] [68]), 
         .C(n33952), .Z(n8_adj_8606)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_68_i8_3_lut.init = 16'hcaca;
    LUT4 i11_4_lut_adj_593 (.A(n5), .B(keymem_sboxw[5]), .C(init_state), 
         .D(n10_adj_8607), .Z(muxed_sboxw[5])) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(181[17:28])
    defparam i11_4_lut_adj_593.init = 16'hc5c0;
    LUT4 i2_3_lut_rep_438 (.A(prev_key1_reg[101]), .B(prev_key1_reg[69]), 
         .C(\round_key_gen.trw[5] ), .Z(n33742)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i2_3_lut_rep_438.init = 16'h9696;
    LUT4 i11_4_lut_adj_594 (.A(n5), .B(keymem_sboxw[6]), .C(init_state), 
         .D(n10_adj_8608), .Z(muxed_sboxw[6])) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(181[17:28])
    defparam i11_4_lut_adj_594.init = 16'hc5c0;
    LUT4 round_3__I_0_Mux_68_i5_3_lut (.A(\key_mem[6] [68]), .B(\key_mem[7] [68]), 
         .C(n33952), .Z(n5_adj_8609)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_68_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_68_i4_3_lut (.A(\key_mem[4] [68]), .B(\key_mem[5] [68]), 
         .C(n33952), .Z(n4_adj_8610)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_68_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_92_i2_3_lut (.A(\key_mem[2] [92]), .B(\key_mem[3] [92]), 
         .C(n33952), .Z(n2_adj_8611)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_92_i2_3_lut.init = 16'hcaca;
    LUT4 i5_2_lut_rep_352_4_lut (.A(prev_key1_reg[101]), .B(prev_key1_reg[69]), 
         .C(\round_key_gen.trw[5] ), .D(prev_key1_reg[37]), .Z(n33656)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i5_2_lut_rep_352_4_lut.init = 16'h6996;
    LUT4 round_3__I_0_Mux_68_i2_3_lut (.A(\key_mem[2] [68]), .B(\key_mem[3] [68]), 
         .C(n33952), .Z(n2_adj_8612)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_68_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_68_i1_3_lut (.A(\key_mem[0] [68]), .B(\key_mem[1] [68]), 
         .C(n33952), .Z(n1_adj_8613)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_68_i1_3_lut.init = 16'hcaca;
    LUT4 i11_4_lut_adj_595 (.A(n5), .B(keymem_sboxw[7]), .C(init_state), 
         .D(n10_adj_8614), .Z(muxed_sboxw[7])) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(181[17:28])
    defparam i11_4_lut_adj_595.init = 16'hc5c0;
    LUT4 i2_3_lut_rep_439 (.A(prev_key1_reg[100]), .B(prev_key1_reg[68]), 
         .C(\round_key_gen.trw[4] ), .Z(n33743)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i2_3_lut_rep_439.init = 16'h9696;
    LUT4 i11_4_lut_adj_596 (.A(n5), .B(keymem_sboxw[8]), .C(init_state), 
         .D(n10_adj_8615), .Z(muxed_sboxw[8])) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(181[17:28])
    defparam i11_4_lut_adj_596.init = 16'hc5c0;
    LUT4 round_3__I_0_Mux_92_i1_3_lut (.A(\key_mem[0] [92]), .B(\key_mem[1] [92]), 
         .C(n33952), .Z(n1_adj_8616)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_92_i1_3_lut.init = 16'hcaca;
    LUT4 i11_4_lut_adj_597 (.A(n5), .B(keymem_sboxw[9]), .C(init_state), 
         .D(n10_adj_8617), .Z(muxed_sboxw[9])) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(181[17:28])
    defparam i11_4_lut_adj_597.init = 16'hc5c0;
    LUT4 round_3__I_0_Mux_67_i11_3_lut (.A(\key_mem[12] [67]), .B(\key_mem[13] [67]), 
         .C(n33952), .Z(n11_adj_39)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_67_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_67_i9_3_lut (.A(\key_mem[10] [67]), .B(\key_mem[11] [67]), 
         .C(n33952), .Z(n9_adj_8619)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_67_i9_3_lut.init = 16'hcaca;
    LUT4 i5_2_lut_rep_354_4_lut (.A(prev_key1_reg[100]), .B(prev_key1_reg[68]), 
         .C(\round_key_gen.trw[4] ), .D(prev_key1_reg[36]), .Z(n33658)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i5_2_lut_rep_354_4_lut.init = 16'h6996;
    LUT4 i11_4_lut_adj_598 (.A(n5), .B(keymem_sboxw[10]), .C(init_state), 
         .D(n10_adj_8620), .Z(muxed_sboxw[10])) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(181[17:28])
    defparam i11_4_lut_adj_598.init = 16'hc5c0;
    LUT4 round_3__I_0_Mux_67_i8_3_lut (.A(\key_mem[8] [67]), .B(\key_mem[9] [67]), 
         .C(n33952), .Z(n8_adj_8621)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_67_i8_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_rep_440 (.A(prev_key1_reg[99]), .B(prev_key1_reg[67]), 
         .C(\round_key_gen.trw[3] ), .Z(n33744)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i2_3_lut_rep_440.init = 16'h9696;
    LUT4 i11_4_lut_adj_599 (.A(n5), .B(keymem_sboxw[11]), .C(init_state), 
         .D(n10_adj_8622), .Z(muxed_sboxw[11])) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(181[17:28])
    defparam i11_4_lut_adj_599.init = 16'hc5c0;
    LUT4 round_3__I_0_Mux_67_i5_3_lut (.A(\key_mem[6] [67]), .B(\key_mem[7] [67]), 
         .C(n33952), .Z(n5_adj_8623)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_67_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_67_i4_3_lut (.A(\key_mem[4] [67]), .B(\key_mem[5] [67]), 
         .C(n33952), .Z(n4_adj_8624)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_67_i4_3_lut.init = 16'hcaca;
    LUT4 i11_4_lut_adj_600 (.A(n5), .B(keymem_sboxw[12]), .C(init_state), 
         .D(n10_adj_8625), .Z(muxed_sboxw[12])) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(181[17:28])
    defparam i11_4_lut_adj_600.init = 16'hc5c0;
    LUT4 i5_2_lut_rep_356_4_lut (.A(prev_key1_reg[99]), .B(prev_key1_reg[67]), 
         .C(\round_key_gen.trw[3] ), .D(prev_key1_reg[35]), .Z(n33660)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i5_2_lut_rep_356_4_lut.init = 16'h6996;
    LUT4 round_3__I_0_Mux_91_i11_3_lut (.A(\key_mem[12] [91]), .B(\key_mem[13] [91]), 
         .C(n33952), .Z(n11_adj_40)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_91_i11_3_lut.init = 16'hcaca;
    LUT4 i11_4_lut_adj_601 (.A(n5), .B(keymem_sboxw[13]), .C(init_state), 
         .D(n10_adj_8627), .Z(muxed_sboxw[13])) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(181[17:28])
    defparam i11_4_lut_adj_601.init = 16'hc5c0;
    LUT4 round_3__I_0_Mux_67_i2_3_lut (.A(\key_mem[2] [67]), .B(\key_mem[3] [67]), 
         .C(n33952), .Z(n2_adj_8628)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_67_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_67_i1_3_lut (.A(\key_mem[0] [67]), .B(\key_mem[1] [67]), 
         .C(n33952), .Z(n1_adj_8629)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_67_i1_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_rep_441 (.A(prev_key1_reg[98]), .B(prev_key1_reg[66]), 
         .C(\round_key_gen.trw[2] ), .Z(n33745)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i2_3_lut_rep_441.init = 16'h9696;
    LUT4 i15019_2_lut_4_lut (.A(\key_reg[5] [16]), .B(n33635), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[80])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15019_2_lut_4_lut.init = 16'hca00;
    LUT4 round_3__I_0_Mux_66_i11_3_lut (.A(\key_mem[12] [66]), .B(\key_mem[13] [66]), 
         .C(n33952), .Z(n11_adj_41)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_66_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_66_i9_3_lut (.A(\key_mem[10] [66]), .B(\key_mem[11] [66]), 
         .C(n33952), .Z(n9_adj_8631)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_66_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_66_i8_3_lut (.A(\key_mem[8] [66]), .B(\key_mem[9] [66]), 
         .C(n33952), .Z(n8_adj_8632)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_66_i8_3_lut.init = 16'hcaca;
    LUT4 i11_4_lut_adj_602 (.A(n5), .B(keymem_sboxw[14]), .C(init_state), 
         .D(n10_adj_8633), .Z(muxed_sboxw[14])) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(181[17:28])
    defparam i11_4_lut_adj_602.init = 16'hc5c0;
    LUT4 round_3__I_0_Mux_66_i5_3_lut (.A(\key_mem[6] [66]), .B(\key_mem[7] [66]), 
         .C(n33952), .Z(n5_adj_8634)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_66_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_66_i4_3_lut (.A(\key_mem[4] [66]), .B(\key_mem[5] [66]), 
         .C(n33952), .Z(n4_adj_8635)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_66_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_91_i9_3_lut (.A(\key_mem[10] [91]), .B(\key_mem[11] [91]), 
         .C(n33952), .Z(n9_adj_8636)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_91_i9_3_lut.init = 16'hcaca;
    LUT4 i11_4_lut_adj_603 (.A(n5), .B(keymem_sboxw[15]), .C(init_state), 
         .D(n10_adj_8637), .Z(muxed_sboxw[15])) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(181[17:28])
    defparam i11_4_lut_adj_603.init = 16'hc5c0;
    LUT4 round_3__I_0_Mux_66_i2_3_lut (.A(\key_mem[2] [66]), .B(\key_mem[3] [66]), 
         .C(n33952), .Z(n2_adj_8638)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_66_i2_3_lut.init = 16'hcaca;
    LUT4 i5_2_lut_rep_358_4_lut (.A(prev_key1_reg[98]), .B(prev_key1_reg[66]), 
         .C(\round_key_gen.trw[2] ), .D(prev_key1_reg[34]), .Z(n33662)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i5_2_lut_rep_358_4_lut.init = 16'h6996;
    LUT4 i11_4_lut_adj_604 (.A(n5), .B(keymem_sboxw[16]), .C(init_state), 
         .D(n10_adj_8639), .Z(\muxed_sboxw[16] )) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(181[17:28])
    defparam i11_4_lut_adj_604.init = 16'hc5c0;
    LUT4 i2_3_lut_rep_442 (.A(prev_key1_reg[97]), .B(prev_key1_reg[65]), 
         .C(\round_key_gen.trw[1] ), .Z(n33746)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i2_3_lut_rep_442.init = 16'h9696;
    LUT4 i11_4_lut_adj_605 (.A(n5), .B(keymem_sboxw[17]), .C(init_state), 
         .D(n10_adj_8640), .Z(\muxed_sboxw[17] )) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(181[17:28])
    defparam i11_4_lut_adj_605.init = 16'hc5c0;
    LUT4 round_3__I_0_Mux_91_i8_3_lut (.A(\key_mem[8] [91]), .B(\key_mem[9] [91]), 
         .C(n33952), .Z(n8_adj_8641)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_91_i8_3_lut.init = 16'hcaca;
    LUT4 i11_4_lut_adj_606 (.A(n5), .B(keymem_sboxw[18]), .C(init_state), 
         .D(n10_adj_8642), .Z(\muxed_sboxw[18] )) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(181[17:28])
    defparam i11_4_lut_adj_606.init = 16'hc5c0;
    LUT4 round_3__I_0_Mux_66_i1_3_lut (.A(\key_mem[0] [66]), .B(\key_mem[1] [66]), 
         .C(n33952), .Z(n1_adj_8643)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_66_i1_3_lut.init = 16'hcaca;
    LUT4 i5_2_lut_rep_360_4_lut (.A(prev_key1_reg[97]), .B(prev_key1_reg[65]), 
         .C(\round_key_gen.trw[1] ), .D(prev_key1_reg[33]), .Z(n33664)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i5_2_lut_rep_360_4_lut.init = 16'h6996;
    LUT4 i2_2_lut_rep_353 (.A(prev_key0_reg[69]), .B(n4_adj_8336), .Z(n33657)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i2_2_lut_rep_353.init = 16'h6666;
    LUT4 i11_4_lut_adj_607 (.A(n5), .B(keymem_sboxw[19]), .C(init_state), 
         .D(n10_adj_8644), .Z(\muxed_sboxw[19] )) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(181[17:28])
    defparam i11_4_lut_adj_607.init = 16'hc5c0;
    LUT4 i2_3_lut_rep_443 (.A(prev_key1_reg[96]), .B(prev_key1_reg[64]), 
         .C(\round_key_gen.trw[0] ), .Z(n33747)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i2_3_lut_rep_443.init = 16'h9696;
    ROM256X1A sboxw_31__I_0_Mux_0 (.AD0(muxed_sboxw[24]), .AD1(muxed_sboxw[25]), 
            .AD2(muxed_sboxw[26]), .AD3(muxed_sboxw[27]), .AD4(muxed_sboxw[28]), 
            .AD5(muxed_sboxw[29]), .AD6(muxed_sboxw[30]), .AD7(muxed_sboxw[31]), 
            .DO0(\round_key_gen.trw[0] )) /* synthesis initstate=0x4F1EAD396F247A0410BDB210C006EAB568AB4BFA8ACB7A13B14EDE67096C6EED */ ;
    defparam sboxw_31__I_0_Mux_0.initval = 256'h4F1EAD396F247A0410BDB210C006EAB568AB4BFA8ACB7A13B14EDE67096C6EED;
    ROM256X1A sboxw_31__I_0_Mux_1 (.AD0(muxed_sboxw[24]), .AD1(muxed_sboxw[25]), 
            .AD2(muxed_sboxw[26]), .AD3(muxed_sboxw[27]), .AD4(muxed_sboxw[28]), 
            .AD5(muxed_sboxw[29]), .AD6(muxed_sboxw[30]), .AD7(muxed_sboxw[31]), 
            .DO0(\round_key_gen.trw[1] )) /* synthesis initstate=0xC870974094EAD8A96A450B2EF33486B4E61A4C5E97816F7A7BAE007D4C53FC7D */ ;
    defparam sboxw_31__I_0_Mux_1.initval = 256'hC870974094EAD8A96A450B2EF33486B4E61A4C5E97816F7A7BAE007D4C53FC7D;
    ROM256X1A sboxw_31__I_0_Mux_4 (.AD0(muxed_sboxw[24]), .AD1(muxed_sboxw[25]), 
            .AD2(muxed_sboxw[26]), .AD3(muxed_sboxw[27]), .AD4(muxed_sboxw[28]), 
            .AD5(muxed_sboxw[29]), .AD6(muxed_sboxw[30]), .AD7(muxed_sboxw[31]), 
            .DO0(\round_key_gen.trw[4] )) /* synthesis initstate=0xF210A3AECE472E532624B286BC48ECB4F7F17A494CE30F58C2B0F97752B8B11E */ ;
    defparam sboxw_31__I_0_Mux_4.initval = 256'hF210A3AECE472E532624B286BC48ECB4F7F17A494CE30F58C2B0F97752B8B11E;
    ROM256X1A sboxw_31__I_0_Mux_2 (.AD0(muxed_sboxw[24]), .AD1(muxed_sboxw[25]), 
            .AD2(muxed_sboxw[26]), .AD3(muxed_sboxw[27]), .AD4(muxed_sboxw[28]), 
            .AD5(muxed_sboxw[29]), .AD6(muxed_sboxw[30]), .AD7(muxed_sboxw[31]), 
            .DO0(\round_key_gen.trw[2] )) /* synthesis initstate=0xAC39B6C0D6CE2EFC577D64E03B0C3FFB23A869A2A428C424A16387FB3B48B4C6 */ ;
    defparam sboxw_31__I_0_Mux_2.initval = 256'hAC39B6C0D6CE2EFC577D64E03B0C3FFB23A869A2A428C424A16387FB3B48B4C6;
    ROM256X1A sboxw_31__I_0_Mux_3 (.AD0(muxed_sboxw[24]), .AD1(muxed_sboxw[25]), 
            .AD2(muxed_sboxw[26]), .AD3(muxed_sboxw[27]), .AD4(muxed_sboxw[28]), 
            .AD5(muxed_sboxw[29]), .AD6(muxed_sboxw[30]), .AD7(muxed_sboxw[31]), 
            .DO0(\round_key_gen.trw[3] )) /* synthesis initstate=0x4E9DDB76C892FB1BE9DA849CF6AC6C1B2568EA2EFFA8527D109020A2193D586A */ ;
    defparam sboxw_31__I_0_Mux_3.initval = 256'h4E9DDB76C892FB1BE9DA849CF6AC6C1B2568EA2EFFA8527D109020A2193D586A;
    ROM256X1A sboxw_31__I_0_Mux_5 (.AD0(muxed_sboxw[24]), .AD1(muxed_sboxw[25]), 
            .AD2(muxed_sboxw[26]), .AD3(muxed_sboxw[27]), .AD4(muxed_sboxw[28]), 
            .AD5(muxed_sboxw[29]), .AD6(muxed_sboxw[30]), .AD7(muxed_sboxw[31]), 
            .DO0(\round_key_gen.trw[5] )) /* synthesis initstate=0x54B248130B4F256F7D8DCC4706319E086BC2AA4E0D787AA4F8045F7B6D98DD7F */ ;
    defparam sboxw_31__I_0_Mux_5.initval = 256'h54B248130B4F256F7D8DCC4706319E086BC2AA4E0D787AA4F8045F7B6D98DD7F;
    ROM256X1A sboxw_31__I_0_Mux_6 (.AD0(muxed_sboxw[24]), .AD1(muxed_sboxw[25]), 
            .AD2(muxed_sboxw[26]), .AD3(muxed_sboxw[27]), .AD4(muxed_sboxw[28]), 
            .AD5(muxed_sboxw[29]), .AD6(muxed_sboxw[30]), .AD7(muxed_sboxw[31]), 
            .DO0(\round_key_gen.trw[6] )) /* synthesis initstate=0x21E0B833255917823F6BCB91B30DB559E4851B3BF3AB2560980A3CC2C2FDB4FF */ ;
    defparam sboxw_31__I_0_Mux_6.initval = 256'h21E0B833255917823F6BCB91B30DB559E4851B3BF3AB2560980A3CC2C2FDB4FF;
    ROM256X1A sboxw_31__I_0_Mux_7 (.AD0(muxed_sboxw[24]), .AD1(muxed_sboxw[25]), 
            .AD2(muxed_sboxw[26]), .AD3(muxed_sboxw[27]), .AD4(muxed_sboxw[28]), 
            .AD5(muxed_sboxw[29]), .AD6(muxed_sboxw[30]), .AD7(muxed_sboxw[31]), 
            .DO0(\round_key_gen.trw[7] )) /* synthesis initstate=0x52379DE7B844E3E14CB3770196CA0329E7BAC28F866AAC825CAA2EC7BF977090 */ ;
    defparam sboxw_31__I_0_Mux_7.initval = 256'h52379DE7B844E3E14CB3770196CA0329E7BAC28F866AAC825CAA2EC7BF977090;
    ROM256X1A sboxw_7__I_0_Mux_0 (.AD0(muxed_sboxw[0]), .AD1(muxed_sboxw[1]), 
            .AD2(muxed_sboxw[2]), .AD3(muxed_sboxw[3]), .AD4(muxed_sboxw[4]), 
            .AD5(muxed_sboxw[5]), .AD6(muxed_sboxw[6]), .AD7(muxed_sboxw[7]), 
            .DO0(\round_key_gen.trw[8] )) /* synthesis initstate=0x4F1EAD396F247A0410BDB210C006EAB568AB4BFA8ACB7A13B14EDE67096C6EED */ ;
    defparam sboxw_7__I_0_Mux_0.initval = 256'h4F1EAD396F247A0410BDB210C006EAB568AB4BFA8ACB7A13B14EDE67096C6EED;
    ROM256X1A sboxw_15__I_0_Mux_0 (.AD0(muxed_sboxw[8]), .AD1(muxed_sboxw[9]), 
            .AD2(muxed_sboxw[10]), .AD3(muxed_sboxw[11]), .AD4(muxed_sboxw[12]), 
            .AD5(muxed_sboxw[13]), .AD6(muxed_sboxw[14]), .AD7(muxed_sboxw[15]), 
            .DO0(\round_key_gen.trw[16] )) /* synthesis initstate=0x4F1EAD396F247A0410BDB210C006EAB568AB4BFA8ACB7A13B14EDE67096C6EED */ ;
    defparam sboxw_15__I_0_Mux_0.initval = 256'h4F1EAD396F247A0410BDB210C006EAB568AB4BFA8ACB7A13B14EDE67096C6EED;
    ROM256X1A sboxw_15__I_0_Mux_7 (.AD0(muxed_sboxw[8]), .AD1(muxed_sboxw[9]), 
            .AD2(muxed_sboxw[10]), .AD3(muxed_sboxw[11]), .AD4(muxed_sboxw[12]), 
            .AD5(muxed_sboxw[13]), .AD6(muxed_sboxw[14]), .AD7(muxed_sboxw[15]), 
            .DO0(\round_key_gen.trw[23] )) /* synthesis initstate=0x52379DE7B844E3E14CB3770196CA0329E7BAC28F866AAC825CAA2EC7BF977090 */ ;
    defparam sboxw_15__I_0_Mux_7.initval = 256'h52379DE7B844E3E14CB3770196CA0329E7BAC28F866AAC825CAA2EC7BF977090;
    ROM256X1A sboxw_15__I_0_Mux_1 (.AD0(muxed_sboxw[8]), .AD1(muxed_sboxw[9]), 
            .AD2(muxed_sboxw[10]), .AD3(muxed_sboxw[11]), .AD4(muxed_sboxw[12]), 
            .AD5(muxed_sboxw[13]), .AD6(muxed_sboxw[14]), .AD7(muxed_sboxw[15]), 
            .DO0(\round_key_gen.trw[17] )) /* synthesis initstate=0xC870974094EAD8A96A450B2EF33486B4E61A4C5E97816F7A7BAE007D4C53FC7D */ ;
    defparam sboxw_15__I_0_Mux_1.initval = 256'hC870974094EAD8A96A450B2EF33486B4E61A4C5E97816F7A7BAE007D4C53FC7D;
    ROM256X1A sboxw_15__I_0_Mux_2 (.AD0(muxed_sboxw[8]), .AD1(muxed_sboxw[9]), 
            .AD2(muxed_sboxw[10]), .AD3(muxed_sboxw[11]), .AD4(muxed_sboxw[12]), 
            .AD5(muxed_sboxw[13]), .AD6(muxed_sboxw[14]), .AD7(muxed_sboxw[15]), 
            .DO0(\round_key_gen.trw[18] )) /* synthesis initstate=0xAC39B6C0D6CE2EFC577D64E03B0C3FFB23A869A2A428C424A16387FB3B48B4C6 */ ;
    defparam sboxw_15__I_0_Mux_2.initval = 256'hAC39B6C0D6CE2EFC577D64E03B0C3FFB23A869A2A428C424A16387FB3B48B4C6;
    ROM256X1A sboxw_7__I_0_Mux_1 (.AD0(muxed_sboxw[0]), .AD1(muxed_sboxw[1]), 
            .AD2(muxed_sboxw[2]), .AD3(muxed_sboxw[3]), .AD4(muxed_sboxw[4]), 
            .AD5(muxed_sboxw[5]), .AD6(muxed_sboxw[6]), .AD7(muxed_sboxw[7]), 
            .DO0(\round_key_gen.trw[9] )) /* synthesis initstate=0xC870974094EAD8A96A450B2EF33486B4E61A4C5E97816F7A7BAE007D4C53FC7D */ ;
    defparam sboxw_7__I_0_Mux_1.initval = 256'hC870974094EAD8A96A450B2EF33486B4E61A4C5E97816F7A7BAE007D4C53FC7D;
    ROM256X1A sboxw_7__I_0_Mux_2 (.AD0(muxed_sboxw[0]), .AD1(muxed_sboxw[1]), 
            .AD2(muxed_sboxw[2]), .AD3(muxed_sboxw[3]), .AD4(muxed_sboxw[4]), 
            .AD5(muxed_sboxw[5]), .AD6(muxed_sboxw[6]), .AD7(muxed_sboxw[7]), 
            .DO0(\round_key_gen.trw[10] )) /* synthesis initstate=0xAC39B6C0D6CE2EFC577D64E03B0C3FFB23A869A2A428C424A16387FB3B48B4C6 */ ;
    defparam sboxw_7__I_0_Mux_2.initval = 256'hAC39B6C0D6CE2EFC577D64E03B0C3FFB23A869A2A428C424A16387FB3B48B4C6;
    ROM256X1A sboxw_7__I_0_Mux_3 (.AD0(muxed_sboxw[0]), .AD1(muxed_sboxw[1]), 
            .AD2(muxed_sboxw[2]), .AD3(muxed_sboxw[3]), .AD4(muxed_sboxw[4]), 
            .AD5(muxed_sboxw[5]), .AD6(muxed_sboxw[6]), .AD7(muxed_sboxw[7]), 
            .DO0(\round_key_gen.trw[11] )) /* synthesis initstate=0x4E9DDB76C892FB1BE9DA849CF6AC6C1B2568EA2EFFA8527D109020A2193D586A */ ;
    defparam sboxw_7__I_0_Mux_3.initval = 256'h4E9DDB76C892FB1BE9DA849CF6AC6C1B2568EA2EFFA8527D109020A2193D586A;
    ROM256X1A sboxw_7__I_0_Mux_4 (.AD0(muxed_sboxw[0]), .AD1(muxed_sboxw[1]), 
            .AD2(muxed_sboxw[2]), .AD3(muxed_sboxw[3]), .AD4(muxed_sboxw[4]), 
            .AD5(muxed_sboxw[5]), .AD6(muxed_sboxw[6]), .AD7(muxed_sboxw[7]), 
            .DO0(\round_key_gen.trw[12] )) /* synthesis initstate=0xF210A3AECE472E532624B286BC48ECB4F7F17A494CE30F58C2B0F97752B8B11E */ ;
    defparam sboxw_7__I_0_Mux_4.initval = 256'hF210A3AECE472E532624B286BC48ECB4F7F17A494CE30F58C2B0F97752B8B11E;
    ROM256X1A sboxw_15__I_0_Mux_3 (.AD0(muxed_sboxw[8]), .AD1(muxed_sboxw[9]), 
            .AD2(muxed_sboxw[10]), .AD3(muxed_sboxw[11]), .AD4(muxed_sboxw[12]), 
            .AD5(muxed_sboxw[13]), .AD6(muxed_sboxw[14]), .AD7(muxed_sboxw[15]), 
            .DO0(\round_key_gen.trw[19] )) /* synthesis initstate=0x4E9DDB76C892FB1BE9DA849CF6AC6C1B2568EA2EFFA8527D109020A2193D586A */ ;
    defparam sboxw_15__I_0_Mux_3.initval = 256'h4E9DDB76C892FB1BE9DA849CF6AC6C1B2568EA2EFFA8527D109020A2193D586A;
    ROM256X1A sboxw_15__I_0_Mux_4 (.AD0(muxed_sboxw[8]), .AD1(muxed_sboxw[9]), 
            .AD2(muxed_sboxw[10]), .AD3(muxed_sboxw[11]), .AD4(muxed_sboxw[12]), 
            .AD5(muxed_sboxw[13]), .AD6(muxed_sboxw[14]), .AD7(muxed_sboxw[15]), 
            .DO0(\round_key_gen.trw[20] )) /* synthesis initstate=0xF210A3AECE472E532624B286BC48ECB4F7F17A494CE30F58C2B0F97752B8B11E */ ;
    defparam sboxw_15__I_0_Mux_4.initval = 256'hF210A3AECE472E532624B286BC48ECB4F7F17A494CE30F58C2B0F97752B8B11E;
    ROM256X1A sboxw_7__I_0_Mux_5 (.AD0(muxed_sboxw[0]), .AD1(muxed_sboxw[1]), 
            .AD2(muxed_sboxw[2]), .AD3(muxed_sboxw[3]), .AD4(muxed_sboxw[4]), 
            .AD5(muxed_sboxw[5]), .AD6(muxed_sboxw[6]), .AD7(muxed_sboxw[7]), 
            .DO0(\round_key_gen.trw[13] )) /* synthesis initstate=0x54B248130B4F256F7D8DCC4706319E086BC2AA4E0D787AA4F8045F7B6D98DD7F */ ;
    defparam sboxw_7__I_0_Mux_5.initval = 256'h54B248130B4F256F7D8DCC4706319E086BC2AA4E0D787AA4F8045F7B6D98DD7F;
    ROM256X1A sboxw_15__I_0_Mux_5 (.AD0(muxed_sboxw[8]), .AD1(muxed_sboxw[9]), 
            .AD2(muxed_sboxw[10]), .AD3(muxed_sboxw[11]), .AD4(muxed_sboxw[12]), 
            .AD5(muxed_sboxw[13]), .AD6(muxed_sboxw[14]), .AD7(muxed_sboxw[15]), 
            .DO0(\round_key_gen.trw[21] )) /* synthesis initstate=0x54B248130B4F256F7D8DCC4706319E086BC2AA4E0D787AA4F8045F7B6D98DD7F */ ;
    defparam sboxw_15__I_0_Mux_5.initval = 256'h54B248130B4F256F7D8DCC4706319E086BC2AA4E0D787AA4F8045F7B6D98DD7F;
    ROM256X1A sboxw_15__I_0_Mux_6 (.AD0(muxed_sboxw[8]), .AD1(muxed_sboxw[9]), 
            .AD2(muxed_sboxw[10]), .AD3(muxed_sboxw[11]), .AD4(muxed_sboxw[12]), 
            .AD5(muxed_sboxw[13]), .AD6(muxed_sboxw[14]), .AD7(muxed_sboxw[15]), 
            .DO0(\round_key_gen.trw[22] )) /* synthesis initstate=0x21E0B833255917823F6BCB91B30DB559E4851B3BF3AB2560980A3CC2C2FDB4FF */ ;
    defparam sboxw_15__I_0_Mux_6.initval = 256'h21E0B833255917823F6BCB91B30DB559E4851B3BF3AB2560980A3CC2C2FDB4FF;
    ROM256X1A sboxw_7__I_0_Mux_6 (.AD0(muxed_sboxw[0]), .AD1(muxed_sboxw[1]), 
            .AD2(muxed_sboxw[2]), .AD3(muxed_sboxw[3]), .AD4(muxed_sboxw[4]), 
            .AD5(muxed_sboxw[5]), .AD6(muxed_sboxw[6]), .AD7(muxed_sboxw[7]), 
            .DO0(\round_key_gen.trw[14] )) /* synthesis initstate=0x21E0B833255917823F6BCB91B30DB559E4851B3BF3AB2560980A3CC2C2FDB4FF */ ;
    defparam sboxw_7__I_0_Mux_6.initval = 256'h21E0B833255917823F6BCB91B30DB559E4851B3BF3AB2560980A3CC2C2FDB4FF;
    ROM256X1A sboxw_7__I_0_Mux_7 (.AD0(muxed_sboxw[0]), .AD1(muxed_sboxw[1]), 
            .AD2(muxed_sboxw[2]), .AD3(muxed_sboxw[3]), .AD4(muxed_sboxw[4]), 
            .AD5(muxed_sboxw[5]), .AD6(muxed_sboxw[6]), .AD7(muxed_sboxw[7]), 
            .DO0(\round_key_gen.trw[15] )) /* synthesis initstate=0x52379DE7B844E3E14CB3770196CA0329E7BAC28F866AAC825CAA2EC7BF977090 */ ;
    defparam sboxw_7__I_0_Mux_7.initval = 256'h52379DE7B844E3E14CB3770196CA0329E7BAC28F866AAC825CAA2EC7BF977090;
    LUT4 i11_4_lut_adj_608 (.A(n5), .B(keymem_sboxw[20]), .C(init_state), 
         .D(n10_adj_8645), .Z(\muxed_sboxw[20] )) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(181[17:28])
    defparam i11_4_lut_adj_608.init = 16'hc5c0;
    LUT4 i5_2_lut_rep_363_4_lut (.A(prev_key1_reg[96]), .B(prev_key1_reg[64]), 
         .C(\round_key_gen.trw[0] ), .D(prev_key1_reg[32]), .Z(n33667)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i5_2_lut_rep_363_4_lut.init = 16'h6996;
    LUT4 round_3__I_0_Mux_91_i5_3_lut (.A(\key_mem[6] [91]), .B(\key_mem[7] [91]), 
         .C(n33952), .Z(n5_adj_8646)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_91_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_65_i11_3_lut (.A(\key_mem[12] [65]), .B(\key_mem[13] [65]), 
         .C(n33952), .Z(n11_adj_42)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_65_i11_3_lut.init = 16'hcaca;
    LUT4 i11_4_lut_adj_609 (.A(n5), .B(keymem_sboxw[21]), .C(init_state), 
         .D(n10_adj_8648), .Z(\muxed_sboxw[21] )) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(181[17:28])
    defparam i11_4_lut_adj_609.init = 16'hc5c0;
    LUT4 round_3__I_0_Mux_91_i4_3_lut (.A(\key_mem[4] [91]), .B(\key_mem[5] [91]), 
         .C(n33952), .Z(n4_adj_8649)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_91_i4_3_lut.init = 16'hcaca;
    LUT4 i11_4_lut_adj_610 (.A(n5), .B(keymem_sboxw[22]), .C(init_state), 
         .D(n10_adj_8650), .Z(\muxed_sboxw[22] )) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(181[17:28])
    defparam i11_4_lut_adj_610.init = 16'hc5c0;
    LUT4 i11_4_lut_adj_611 (.A(n5), .B(keymem_sboxw[23]), .C(init_state), 
         .D(n10_adj_8651), .Z(\muxed_sboxw[23] )) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(181[17:28])
    defparam i11_4_lut_adj_611.init = 16'hc5c0;
    LUT4 round_3__I_0_Mux_65_i9_3_lut (.A(\key_mem[10] [65]), .B(\key_mem[11] [65]), 
         .C(n33952), .Z(n9_adj_8652)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_65_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_65_i8_3_lut (.A(\key_mem[8] [65]), .B(\key_mem[9] [65]), 
         .C(n33952), .Z(n8_adj_8653)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_65_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_65_i5_3_lut (.A(\key_mem[6] [65]), .B(\key_mem[7] [65]), 
         .C(n33952), .Z(n5_adj_8654)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_65_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_65_i4_3_lut (.A(\key_mem[4] [65]), .B(\key_mem[5] [65]), 
         .C(n33952), .Z(n4_adj_8655)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_65_i4_3_lut.init = 16'hcaca;
    LUT4 mux_85_i70_3_lut_rep_248_4_lut (.A(prev_key0_reg[69]), .B(n4_adj_8336), 
         .C(n33859), .D(\key_reg[5] [5]), .Z(n33552)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam mux_85_i70_3_lut_rep_248_4_lut.init = 16'h6f60;
    LUT4 round_3__I_0_Mux_65_i2_3_lut (.A(\key_mem[2] [65]), .B(\key_mem[3] [65]), 
         .C(n33952), .Z(n2_adj_8656)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_65_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_65_i1_3_lut (.A(\key_mem[0] [65]), .B(\key_mem[1] [65]), 
         .C(n33952), .Z(n1_adj_8657)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_65_i1_3_lut.init = 16'hcaca;
    FD1S3AX ready_reg_155 (.D(n8478), .CK(clk_c), .Q(key_ready));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam ready_reg_155.GSR = "ENABLED";
    LUT4 i3_4_lut (.A(n2958), .B(n6361[2]), .C(n6361[0]), .D(n33951), 
         .Z(key_mem_ctrl_we)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam i3_4_lut.init = 16'hfffe;
    LUT4 i305_2_lut (.A(n7), .B(n35839), .Z(n2958)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam i305_2_lut.init = 16'h4444;
    LUT4 i15018_2_lut_4_lut (.A(\key_reg[5] [15]), .B(n33637), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[79])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15018_2_lut_4_lut.init = 16'hca00;
    LUT4 i2_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), .C(\key_mem_ctrl.num_rounds[2] ), 
         .D(n33912), .Z(n7)) /* synthesis lut_function=(A (((D)+!C)+!B)+!A ((C+(D))+!B)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(405[17:44])
    defparam i2_4_lut.init = 16'hff7b;
    LUT4 round_3__I_0_Mux_64_i11_3_lut (.A(\key_mem[12] [64]), .B(\key_mem[13] [64]), 
         .C(n33952), .Z(n11_adj_43)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_64_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_42_i11_3_lut (.A(\key_mem[12] [42]), .B(\key_mem[13] [42]), 
         .C(n33952), .Z(n11_adj_44)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_42_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_64_i9_3_lut (.A(\key_mem[10] [64]), .B(\key_mem[11] [64]), 
         .C(n33952), .Z(n9_adj_8660)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_64_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_42_i9_3_lut (.A(\key_mem[10] [42]), .B(\key_mem[11] [42]), 
         .C(n33952), .Z(n9_adj_8661)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_42_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_64_i8_3_lut (.A(\key_mem[8] [64]), .B(\key_mem[9] [64]), 
         .C(n33952), .Z(n8_adj_8662)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_64_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_42_i8_3_lut (.A(\key_mem[8] [42]), .B(\key_mem[9] [42]), 
         .C(n33952), .Z(n8_adj_8663)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_42_i8_3_lut.init = 16'hcaca;
    FD1P3AX key_mem_ctrl_reg_FSM_i0_i0 (.D(n2958), .SP(key_mem_ctrl_we), 
            .CK(clk_c), .Q(n6361[0]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam key_mem_ctrl_reg_FSM_i0_i0.GSR = "ENABLED";
    LUT4 round_3__I_0_Mux_64_i5_3_lut (.A(\key_mem[6] [64]), .B(\key_mem[7] [64]), 
         .C(n33952), .Z(n5_adj_8664)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_64_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_64_i4_3_lut (.A(\key_mem[4] [64]), .B(\key_mem[5] [64]), 
         .C(n33952), .Z(n4_adj_8665)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_64_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_42_i5_3_lut (.A(\key_mem[6] [42]), .B(\key_mem[7] [42]), 
         .C(n33952), .Z(n5_adj_8666)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_42_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_64_i2_3_lut (.A(\key_mem[2] [64]), .B(\key_mem[3] [64]), 
         .C(n33952), .Z(n2_adj_8667)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_64_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_42_i4_3_lut (.A(\key_mem[4] [42]), .B(\key_mem[5] [42]), 
         .C(n33952), .Z(n4_adj_8668)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_42_i4_3_lut.init = 16'hcaca;
    LUT4 i15062_2_lut_4_lut (.A(\key_reg[4] [27]), .B(n4_adj_8444), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[123])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15062_2_lut_4_lut.init = 16'hca00;
    LUT4 round_3__I_0_Mux_64_i1_3_lut (.A(\key_mem[0] [64]), .B(\key_mem[1] [64]), 
         .C(n33952), .Z(n1_adj_8669)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_64_i1_3_lut.init = 16'hcaca;
    LUT4 i15017_2_lut_4_lut (.A(\key_reg[5] [14]), .B(n33639), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[78])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15017_2_lut_4_lut.init = 16'hca00;
    LUT4 round_3__I_0_Mux_42_i2_3_lut (.A(\key_mem[2] [42]), .B(\key_mem[3] [42]), 
         .C(n33952), .Z(n2_adj_8670)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_42_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_63_i11_3_lut (.A(\key_mem[12] [63]), .B(\key_mem[13] [63]), 
         .C(n33952), .Z(n11_adj_45)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_63_i11_3_lut.init = 16'hcaca;
    LUT4 i15061_2_lut_4_lut (.A(\key_reg[4] [26]), .B(n4_adj_8438), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[122])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15061_2_lut_4_lut.init = 16'hca00;
    LUT4 round_3__I_0_Mux_63_i9_3_lut (.A(\key_mem[10] [63]), .B(\key_mem[11] [63]), 
         .C(n33952), .Z(n9_adj_8672)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_63_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_63_i8_3_lut (.A(\key_mem[8] [63]), .B(\key_mem[9] [63]), 
         .C(n33952), .Z(n8_adj_8673)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_63_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_42_i1_3_lut (.A(\key_mem[0] [42]), .B(\key_mem[1] [42]), 
         .C(n33952), .Z(n1_adj_8674)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_42_i1_3_lut.init = 16'hcaca;
    LUT4 i15034_2_lut_4_lut (.A(\key_reg[5] [31]), .B(n33558), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[95])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15034_2_lut_4_lut.init = 16'hca00;
    LUT4 round_3__I_0_Mux_91_i2_3_lut (.A(\key_mem[2] [91]), .B(\key_mem[3] [91]), 
         .C(n33952), .Z(n2_adj_8675)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_91_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_91_i1_3_lut (.A(\key_mem[0] [91]), .B(\key_mem[1] [91]), 
         .C(n33952), .Z(n1_adj_8676)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_91_i1_3_lut.init = 16'hcaca;
    LUT4 i6_2_lut_3_lut_adj_612 (.A(prev_key1_reg[36]), .B(n33743), .C(keymem_sboxw[4]), 
         .Z(n15597)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;
    defparam i6_2_lut_3_lut_adj_612.init = 16'h9696;
    LUT4 round_3__I_0_Mux_63_i5_3_lut (.A(\key_mem[6] [63]), .B(\key_mem[7] [63]), 
         .C(n33952), .Z(n5_adj_8677)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_63_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_63_i4_3_lut (.A(\key_mem[4] [63]), .B(\key_mem[5] [63]), 
         .C(n33952), .Z(n4_adj_8678)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_63_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_41_i11_3_lut (.A(\key_mem[12] [41]), .B(\key_mem[13] [41]), 
         .C(n33952), .Z(n11_adj_46)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_41_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_63_i2_3_lut (.A(\key_mem[2] [63]), .B(\key_mem[3] [63]), 
         .C(n33952), .Z(n2_adj_8680)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_63_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_41_i9_3_lut (.A(\key_mem[10] [41]), .B(\key_mem[11] [41]), 
         .C(n33952), .Z(n9_adj_8681)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_41_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_41_i8_3_lut (.A(\key_mem[8] [41]), .B(\key_mem[9] [41]), 
         .C(n33952), .Z(n8_adj_8682)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_41_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_63_i1_3_lut (.A(\key_mem[0] [63]), .B(\key_mem[1] [63]), 
         .C(n33952), .Z(n1_adj_8683)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_63_i1_3_lut.init = 16'hcaca;
    LUT4 i15016_2_lut_4_lut (.A(\key_reg[5] [13]), .B(n33641), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[77])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15016_2_lut_4_lut.init = 16'hca00;
    LUT4 i1_2_lut_adj_613 (.A(n35839), .B(reset_n_c), .Z(n28850)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam i1_2_lut_adj_613.init = 16'h8888;
    LUT4 i2_2_lut_rep_355 (.A(prev_key0_reg[68]), .B(n4_adj_8335), .Z(n33659)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i2_2_lut_rep_355.init = 16'h6666;
    LUT4 round_3__I_0_Mux_90_i11_3_lut (.A(\key_mem[12] [90]), .B(\key_mem[13] [90]), 
         .C(n33952), .Z(n11_adj_47)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_90_i11_3_lut.init = 16'hcaca;
    LUT4 mux_85_i69_3_lut_rep_249_4_lut (.A(prev_key0_reg[68]), .B(n4_adj_8335), 
         .C(n33859), .D(\key_reg[5] [4]), .Z(n33553)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam mux_85_i69_3_lut_rep_249_4_lut.init = 16'h6f60;
    LUT4 round_3__I_0_Mux_90_i9_3_lut (.A(\key_mem[10] [90]), .B(\key_mem[11] [90]), 
         .C(n33952), .Z(n9_adj_8685)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_90_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_90_i8_3_lut (.A(\key_mem[8] [90]), .B(\key_mem[9] [90]), 
         .C(n33952), .Z(n8_adj_8686)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_90_i8_3_lut.init = 16'hcaca;
    LUT4 i15060_2_lut_4_lut (.A(\key_reg[4] [25]), .B(n4_adj_8430), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[121])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15060_2_lut_4_lut.init = 16'hca00;
    LUT4 i15059_2_lut_4_lut (.A(\key_reg[4] [24]), .B(n4_adj_8428), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[120])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15059_2_lut_4_lut.init = 16'hca00;
    LUT4 round_3__I_0_Mux_90_i5_3_lut (.A(\key_mem[6] [90]), .B(\key_mem[7] [90]), 
         .C(n33952), .Z(n5_adj_8687)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_90_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_90_i4_3_lut (.A(\key_mem[4] [90]), .B(\key_mem[5] [90]), 
         .C(n33952), .Z(n4_adj_8688)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_90_i4_3_lut.init = 16'hcaca;
    LUT4 i6_2_lut_3_lut_adj_614 (.A(prev_key1_reg[35]), .B(n33744), .C(keymem_sboxw[3]), 
         .Z(n15537)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;
    defparam i6_2_lut_3_lut_adj_614.init = 16'h9696;
    LUT4 i2_2_lut_rep_357 (.A(prev_key0_reg[67]), .B(n4_adj_8333), .Z(n33661)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i2_2_lut_rep_357.init = 16'h6666;
    LUT4 mux_85_i68_3_lut_rep_250_4_lut (.A(prev_key0_reg[67]), .B(n4_adj_8333), 
         .C(n33859), .D(\key_reg[5] [3]), .Z(n33554)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam mux_85_i68_3_lut_rep_250_4_lut.init = 16'h6f60;
    LUT4 i6_2_lut_3_lut_adj_615 (.A(prev_key1_reg[34]), .B(n33745), .C(keymem_sboxw[2]), 
         .Z(n15477)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;
    defparam i6_2_lut_3_lut_adj_615.init = 16'h9696;
    LUT4 i2_2_lut_rep_359 (.A(prev_key0_reg[66]), .B(n4_adj_8332), .Z(n33663)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i2_2_lut_rep_359.init = 16'h6666;
    LUT4 mux_85_i67_3_lut_rep_251_4_lut (.A(prev_key0_reg[66]), .B(n4_adj_8332), 
         .C(n33859), .D(\key_reg[5] [2]), .Z(n33555)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam mux_85_i67_3_lut_rep_251_4_lut.init = 16'h6f60;
    LUT4 round_3__I_0_Mux_90_i2_3_lut (.A(\key_mem[2] [90]), .B(\key_mem[3] [90]), 
         .C(n33952), .Z(n2_adj_8689)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_90_i2_3_lut.init = 16'hcaca;
    LUT4 i15026_2_lut_4_lut (.A(\key_reg[5] [23]), .B(n33621), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[87])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15026_2_lut_4_lut.init = 16'hca00;
    LUT4 i6_2_lut_3_lut_adj_616 (.A(prev_key1_reg[33]), .B(n33746), .C(keymem_sboxw[1]), 
         .Z(n15417)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;
    defparam i6_2_lut_3_lut_adj_616.init = 16'h9696;
    LUT4 round_3__I_0_Mux_90_i1_3_lut (.A(\key_mem[0] [90]), .B(\key_mem[1] [90]), 
         .C(n33952), .Z(n1_adj_8690)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_90_i1_3_lut.init = 16'hcaca;
    LUT4 i2_2_lut_rep_361 (.A(prev_key0_reg[65]), .B(n8929), .Z(n33665)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i2_2_lut_rep_361.init = 16'h6666;
    LUT4 round_3__I_0_Mux_89_i11_3_lut (.A(\key_mem[12] [89]), .B(\key_mem[13] [89]), 
         .C(n33952), .Z(n11_adj_48)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_89_i11_3_lut.init = 16'hcaca;
    LUT4 mux_85_i66_3_lut_rep_252_4_lut (.A(prev_key0_reg[65]), .B(n8929), 
         .C(n33859), .D(\key_reg[5] [1]), .Z(n33556)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam mux_85_i66_3_lut_rep_252_4_lut.init = 16'h6f60;
    LUT4 round_3__I_0_Mux_89_i9_3_lut (.A(\key_mem[10] [89]), .B(\key_mem[11] [89]), 
         .C(n33952), .Z(n9_adj_8692)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_89_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_89_i8_3_lut (.A(\key_mem[8] [89]), .B(\key_mem[9] [89]), 
         .C(n33952), .Z(n8_adj_8693)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_89_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_89_i5_3_lut (.A(\key_mem[6] [89]), .B(\key_mem[7] [89]), 
         .C(n33952), .Z(n5_adj_8694)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_89_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_89_i4_3_lut (.A(\key_mem[4] [89]), .B(\key_mem[5] [89]), 
         .C(n33952), .Z(n4_adj_8695)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_89_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_89_i2_3_lut (.A(\key_mem[2] [89]), .B(\key_mem[3] [89]), 
         .C(n33952), .Z(n2_adj_8696)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_89_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_89_i1_3_lut (.A(\key_mem[0] [89]), .B(\key_mem[1] [89]), 
         .C(n33952), .Z(n1_adj_8697)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_89_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_88_i11_3_lut (.A(\key_mem[12] [88]), .B(\key_mem[13] [88]), 
         .C(n33952), .Z(n11_adj_49)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_88_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_88_i9_3_lut (.A(\key_mem[10] [88]), .B(\key_mem[11] [88]), 
         .C(n33952), .Z(n9_adj_8699)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_88_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_88_i8_3_lut (.A(\key_mem[8] [88]), .B(\key_mem[9] [88]), 
         .C(n33952), .Z(n8_adj_8700)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_88_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_88_i5_3_lut (.A(\key_mem[6] [88]), .B(\key_mem[7] [88]), 
         .C(n33952), .Z(n5_adj_8701)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_88_i5_3_lut.init = 16'hcaca;
    LUT4 i2_2_lut_rep_362 (.A(prev_key0_reg[64]), .B(n8487), .Z(n33666)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i2_2_lut_rep_362.init = 16'h6666;
    LUT4 round_3__I_0_Mux_88_i4_3_lut (.A(\key_mem[4] [88]), .B(\key_mem[5] [88]), 
         .C(n33952), .Z(n4_adj_8702)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_88_i4_3_lut.init = 16'hcaca;
    LUT4 mux_85_i65_3_lut_rep_253_4_lut (.A(prev_key0_reg[64]), .B(n8487), 
         .C(n33859), .D(\key_reg[5] [0]), .Z(n33557)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam mux_85_i65_3_lut_rep_253_4_lut.init = 16'h6f60;
    LUT4 round_3__I_0_Mux_41_i5_3_lut (.A(\key_mem[6] [41]), .B(\key_mem[7] [41]), 
         .C(n33952), .Z(n5_adj_8703)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_41_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_62_i11_3_lut (.A(\key_mem[12] [62]), .B(\key_mem[13] [62]), 
         .C(n33952), .Z(n11_adj_50)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_62_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_41_i4_3_lut (.A(\key_mem[4] [41]), .B(\key_mem[5] [41]), 
         .C(n33952), .Z(n4_adj_8705)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_41_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_41_i2_3_lut (.A(\key_mem[2] [41]), .B(\key_mem[3] [41]), 
         .C(n33952), .Z(n2_adj_8706)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_41_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_62_i9_3_lut (.A(\key_mem[10] [62]), .B(\key_mem[11] [62]), 
         .C(n33952), .Z(n9_adj_8707)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_62_i9_3_lut.init = 16'hcaca;
    PFUMX i25681 (.BLUT(n1_adj_8708), .ALUT(n2_adj_8709), .C0(\muxed_round_nr[1] ), 
          .Z(n30840));
    LUT4 round_3__I_0_Mux_62_i8_3_lut (.A(\key_mem[8] [62]), .B(\key_mem[9] [62]), 
         .C(n33952), .Z(n8_adj_8710)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_62_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_62_i5_3_lut (.A(\key_mem[6] [62]), .B(\key_mem[7] [62]), 
         .C(n33952), .Z(n5_adj_8711)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_62_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_41_i1_3_lut (.A(\key_mem[0] [41]), .B(\key_mem[1] [41]), 
         .C(n33952), .Z(n1_adj_8712)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_41_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_62_i4_3_lut (.A(\key_mem[4] [62]), .B(\key_mem[5] [62]), 
         .C(n33952), .Z(n4_adj_8713)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_62_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_62_i2_3_lut (.A(\key_mem[2] [62]), .B(\key_mem[3] [62]), 
         .C(n33952), .Z(n2_adj_8714)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_62_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_62_i1_3_lut (.A(\key_mem[0] [62]), .B(\key_mem[1] [62]), 
         .C(n33952), .Z(n1_adj_8715)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_62_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_40_i11_3_lut (.A(\key_mem[12] [40]), .B(\key_mem[13] [40]), 
         .C(n33952), .Z(n11_adj_51)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_40_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_40_i9_3_lut (.A(\key_mem[10] [40]), .B(\key_mem[11] [40]), 
         .C(n33952), .Z(n9_adj_8717)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_40_i9_3_lut.init = 16'hcaca;
    LUT4 i15015_2_lut_4_lut (.A(\key_reg[5] [12]), .B(n33643), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[76])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15015_2_lut_4_lut.init = 16'hca00;
    LUT4 round_3__I_0_Mux_40_i8_3_lut (.A(\key_mem[8] [40]), .B(\key_mem[9] [40]), 
         .C(n33952), .Z(n8_adj_8718)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_40_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_40_i5_3_lut (.A(\key_mem[6] [40]), .B(\key_mem[7] [40]), 
         .C(n33952), .Z(n5_adj_8719)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_40_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_40_i4_3_lut (.A(\key_mem[4] [40]), .B(\key_mem[5] [40]), 
         .C(n33952), .Z(n4_adj_8720)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_40_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_61_i11_3_lut (.A(\key_mem[12] [61]), .B(\key_mem[13] [61]), 
         .C(n33952), .Z(n11_adj_52)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_61_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_61_i9_3_lut (.A(\key_mem[10] [61]), .B(\key_mem[11] [61]), 
         .C(n33952), .Z(n9_adj_8722)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_61_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_61_i8_3_lut (.A(\key_mem[8] [61]), .B(\key_mem[9] [61]), 
         .C(n33952), .Z(n8_adj_8723)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_61_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_61_i5_3_lut (.A(\key_mem[6] [61]), .B(\key_mem[7] [61]), 
         .C(n33952), .Z(n5_adj_8724)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_61_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_61_i4_3_lut (.A(\key_mem[4] [61]), .B(\key_mem[5] [61]), 
         .C(n33952), .Z(n4_adj_8725)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_61_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_40_i2_3_lut (.A(\key_mem[2] [40]), .B(\key_mem[3] [40]), 
         .C(n33952), .Z(n2_adj_8726)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_40_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_61_i2_3_lut (.A(\key_mem[2] [61]), .B(\key_mem[3] [61]), 
         .C(n33952), .Z(n2_adj_8727)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_61_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_40_i1_3_lut (.A(\key_mem[0] [40]), .B(\key_mem[1] [40]), 
         .C(n33952), .Z(n1_adj_8728)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_40_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_61_i1_3_lut (.A(\key_mem[0] [61]), .B(\key_mem[1] [61]), 
         .C(n33952), .Z(n1_adj_8729)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_61_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_60_i11_3_lut (.A(\key_mem[12] [60]), .B(\key_mem[13] [60]), 
         .C(n33952), .Z(n11_adj_53)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_60_i11_3_lut.init = 16'hcaca;
    LUT4 i15014_2_lut_4_lut (.A(\key_reg[5] [11]), .B(n33645), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[75])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15014_2_lut_4_lut.init = 16'hca00;
    LUT4 round_3__I_0_Mux_39_i11_3_lut (.A(\key_mem[12] [39]), .B(\key_mem[13] [39]), 
         .C(n33952), .Z(n11_adj_54)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_39_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_60_i9_3_lut (.A(\key_mem[10] [60]), .B(\key_mem[11] [60]), 
         .C(n33952), .Z(n9_adj_8732)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_60_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_39_i9_3_lut (.A(\key_mem[10] [39]), .B(\key_mem[11] [39]), 
         .C(n33952), .Z(n9_adj_8733)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_39_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_60_i8_3_lut (.A(\key_mem[8] [60]), .B(\key_mem[9] [60]), 
         .C(n33952), .Z(n8_adj_8734)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_60_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_39_i8_3_lut (.A(\key_mem[8] [39]), .B(\key_mem[9] [39]), 
         .C(n33952), .Z(n8_adj_8735)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_39_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_60_i5_3_lut (.A(\key_mem[6] [60]), .B(\key_mem[7] [60]), 
         .C(n33952), .Z(n5_adj_8736)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_60_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_39_i5_3_lut (.A(\key_mem[6] [39]), .B(\key_mem[7] [39]), 
         .C(n33952), .Z(n5_adj_8737)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_39_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_60_i4_3_lut (.A(\key_mem[4] [60]), .B(\key_mem[5] [60]), 
         .C(n33952), .Z(n4_adj_8738)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_60_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_39_i4_3_lut (.A(\key_mem[4] [39]), .B(\key_mem[5] [39]), 
         .C(n33952), .Z(n4_adj_8739)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_39_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_39_i2_3_lut (.A(\key_mem[2] [39]), .B(\key_mem[3] [39]), 
         .C(n33952), .Z(n2_adj_8740)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_39_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_39_i1_3_lut (.A(\key_mem[0] [39]), .B(\key_mem[1] [39]), 
         .C(n33952), .Z(n1_adj_8741)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_39_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_60_i2_3_lut (.A(\key_mem[2] [60]), .B(\key_mem[3] [60]), 
         .C(n33952), .Z(n2_adj_8742)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_60_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_60_i1_3_lut (.A(\key_mem[0] [60]), .B(\key_mem[1] [60]), 
         .C(n33952), .Z(n1_adj_8743)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_60_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_38_i11_3_lut (.A(\key_mem[12] [38]), .B(\key_mem[13] [38]), 
         .C(n33952), .Z(n11_adj_55)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_38_i11_3_lut.init = 16'hcaca;
    LUT4 i15013_2_lut_4_lut (.A(\key_reg[5] [10]), .B(n33647), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[74])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15013_2_lut_4_lut.init = 16'hca00;
    LUT4 round_3__I_0_Mux_59_i11_3_lut (.A(\key_mem[12] [59]), .B(\key_mem[13] [59]), 
         .C(n33952), .Z(n11_adj_56)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_59_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_59_i9_3_lut (.A(\key_mem[10] [59]), .B(\key_mem[11] [59]), 
         .C(n33952), .Z(n9_adj_8746)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_59_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_59_i8_3_lut (.A(\key_mem[8] [59]), .B(\key_mem[9] [59]), 
         .C(n33952), .Z(n8_adj_8747)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_59_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_59_i5_3_lut (.A(\key_mem[6] [59]), .B(\key_mem[7] [59]), 
         .C(n33952), .Z(n5_adj_8748)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_59_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_38_i9_3_lut (.A(\key_mem[10] [38]), .B(\key_mem[11] [38]), 
         .C(n33952), .Z(n9_adj_8749)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_38_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_38_i8_3_lut (.A(\key_mem[8] [38]), .B(\key_mem[9] [38]), 
         .C(n33952), .Z(n8_adj_8750)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_38_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_59_i4_3_lut (.A(\key_mem[4] [59]), .B(\key_mem[5] [59]), 
         .C(n33952), .Z(n4_adj_8751)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_59_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_38_i5_3_lut (.A(\key_mem[6] [38]), .B(\key_mem[7] [38]), 
         .C(n33952), .Z(n5_adj_8752)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_38_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_38_i4_3_lut (.A(\key_mem[4] [38]), .B(\key_mem[5] [38]), 
         .C(n33952), .Z(n4_adj_8753)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_38_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_59_i2_3_lut (.A(\key_mem[2] [59]), .B(\key_mem[3] [59]), 
         .C(n33952), .Z(n2_adj_8754)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_59_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_38_i2_3_lut (.A(\key_mem[2] [38]), .B(\key_mem[3] [38]), 
         .C(n33952), .Z(n2_adj_8755)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_38_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_59_i1_3_lut (.A(\key_mem[0] [59]), .B(\key_mem[1] [59]), 
         .C(n33952), .Z(n1_adj_8756)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_59_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_38_i1_3_lut (.A(\key_mem[0] [38]), .B(\key_mem[1] [38]), 
         .C(n33952), .Z(n1_adj_8757)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_38_i1_3_lut.init = 16'hcaca;
    LUT4 i15012_2_lut_4_lut (.A(\key_reg[5] [9]), .B(n33649), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[73])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15012_2_lut_4_lut.init = 16'hca00;
    LUT4 round_3__I_0_Mux_58_i11_3_lut (.A(\key_mem[12] [58]), .B(\key_mem[13] [58]), 
         .C(n33952), .Z(n11_adj_57)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_58_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_58_i9_3_lut (.A(\key_mem[10] [58]), .B(\key_mem[11] [58]), 
         .C(n33952), .Z(n9_adj_8759)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_58_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_58_i8_3_lut (.A(\key_mem[8] [58]), .B(\key_mem[9] [58]), 
         .C(n33952), .Z(n8_adj_8760)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_58_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_37_i11_3_lut (.A(\key_mem[12] [37]), .B(\key_mem[13] [37]), 
         .C(n33952), .Z(n11_adj_58)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_37_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_37_i9_3_lut (.A(\key_mem[10] [37]), .B(\key_mem[11] [37]), 
         .C(n33952), .Z(n9_adj_8762)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_37_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_58_i5_3_lut (.A(\key_mem[6] [58]), .B(\key_mem[7] [58]), 
         .C(n33952), .Z(n5_adj_8763)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_58_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_58_i4_3_lut (.A(\key_mem[4] [58]), .B(\key_mem[5] [58]), 
         .C(n33952), .Z(n4_adj_8764)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_58_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_37_i8_3_lut (.A(\key_mem[8] [37]), .B(\key_mem[9] [37]), 
         .C(n33952), .Z(n8_adj_8765)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_37_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_58_i2_3_lut (.A(\key_mem[2] [58]), .B(\key_mem[3] [58]), 
         .C(n33952), .Z(n2_adj_8766)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_58_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_37_i5_3_lut (.A(\key_mem[6] [37]), .B(\key_mem[7] [37]), 
         .C(n33952), .Z(n5_adj_8767)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_37_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_58_i1_3_lut (.A(\key_mem[0] [58]), .B(\key_mem[1] [58]), 
         .C(n33952), .Z(n1_adj_8768)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_58_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_37_i4_3_lut (.A(\key_mem[4] [37]), .B(\key_mem[5] [37]), 
         .C(n33952), .Z(n4_adj_8769)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_37_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_57_i11_3_lut (.A(\key_mem[12] [57]), .B(\key_mem[13] [57]), 
         .C(n33952), .Z(n11_adj_59)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_57_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_37_i2_3_lut (.A(\key_mem[2] [37]), .B(\key_mem[3] [37]), 
         .C(n33952), .Z(n2_adj_8771)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_37_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_37_i1_3_lut (.A(\key_mem[0] [37]), .B(\key_mem[1] [37]), 
         .C(n33952), .Z(n1_adj_8772)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_37_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_57_i9_3_lut (.A(\key_mem[10] [57]), .B(\key_mem[11] [57]), 
         .C(n33952), .Z(n9_adj_8773)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_57_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_57_i8_3_lut (.A(\key_mem[8] [57]), .B(\key_mem[9] [57]), 
         .C(n33952), .Z(n8_adj_8774)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_57_i8_3_lut.init = 16'hcaca;
    LUT4 i15011_2_lut_4_lut (.A(\key_reg[5] [8]), .B(n33651), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[72])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15011_2_lut_4_lut.init = 16'hca00;
    LUT4 round_3__I_0_Mux_36_i11_3_lut (.A(\key_mem[12] [36]), .B(\key_mem[13] [36]), 
         .C(n33952), .Z(n11_adj_60)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_36_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_57_i5_3_lut (.A(\key_mem[6] [57]), .B(\key_mem[7] [57]), 
         .C(n33952), .Z(n5_adj_8776)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_57_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_57_i4_3_lut (.A(\key_mem[4] [57]), .B(\key_mem[5] [57]), 
         .C(n33952), .Z(n4_adj_8777)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_57_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_57_i2_3_lut (.A(\key_mem[2] [57]), .B(\key_mem[3] [57]), 
         .C(n33952), .Z(n2_adj_8778)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_57_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_57_i1_3_lut (.A(\key_mem[0] [57]), .B(\key_mem[1] [57]), 
         .C(n33952), .Z(n1_adj_8779)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_57_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_36_i9_3_lut (.A(\key_mem[10] [36]), .B(\key_mem[11] [36]), 
         .C(n33952), .Z(n9_adj_8780)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_36_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_36_i8_3_lut (.A(\key_mem[8] [36]), .B(\key_mem[9] [36]), 
         .C(n33952), .Z(n8_adj_8781)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_36_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_36_i5_3_lut (.A(\key_mem[6] [36]), .B(\key_mem[7] [36]), 
         .C(n33952), .Z(n5_adj_8782)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_36_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_36_i4_3_lut (.A(\key_mem[4] [36]), .B(\key_mem[5] [36]), 
         .C(n33952), .Z(n4_adj_8783)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_36_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_56_i11_3_lut (.A(\key_mem[12] [56]), .B(\key_mem[13] [56]), 
         .C(n33952), .Z(n11_adj_61)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_56_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_36_i2_3_lut (.A(\key_mem[2] [36]), .B(\key_mem[3] [36]), 
         .C(n33952), .Z(n2_adj_8785)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_36_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_36_i1_3_lut (.A(\key_mem[0] [36]), .B(\key_mem[1] [36]), 
         .C(n33952), .Z(n1_adj_8786)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_36_i1_3_lut.init = 16'hcaca;
    LUT4 i15010_2_lut_4_lut (.A(\key_reg[5] [7]), .B(n33653), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[71])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15010_2_lut_4_lut.init = 16'hca00;
    LUT4 round_3__I_0_Mux_56_i9_3_lut (.A(\key_mem[10] [56]), .B(\key_mem[11] [56]), 
         .C(n33952), .Z(n9_adj_8787)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_56_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_56_i8_3_lut (.A(\key_mem[8] [56]), .B(\key_mem[9] [56]), 
         .C(n33952), .Z(n8_adj_8788)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_56_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_56_i5_3_lut (.A(\key_mem[6] [56]), .B(\key_mem[7] [56]), 
         .C(n33952), .Z(n5_adj_8789)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_56_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_35_i11_3_lut (.A(\key_mem[12] [35]), .B(\key_mem[13] [35]), 
         .C(n33952), .Z(n11_adj_62)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_35_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_56_i4_3_lut (.A(\key_mem[4] [56]), .B(\key_mem[5] [56]), 
         .C(n33952), .Z(n4_adj_8791)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_56_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_56_i2_3_lut (.A(\key_mem[2] [56]), .B(\key_mem[3] [56]), 
         .C(n33952), .Z(n2_adj_8792)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_56_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_56_i1_3_lut (.A(\key_mem[0] [56]), .B(\key_mem[1] [56]), 
         .C(n33952), .Z(n1_adj_8793)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_56_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_35_i9_3_lut (.A(\key_mem[10] [35]), .B(\key_mem[11] [35]), 
         .C(n33952), .Z(n9_adj_8794)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_35_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_35_i8_3_lut (.A(\key_mem[8] [35]), .B(\key_mem[9] [35]), 
         .C(n33952), .Z(n8_adj_8795)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_35_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_55_i11_3_lut (.A(\key_mem[12] [55]), .B(\key_mem[13] [55]), 
         .C(n33952), .Z(n11_adj_63)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_55_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_55_i9_3_lut (.A(\key_mem[10] [55]), .B(\key_mem[11] [55]), 
         .C(n33952), .Z(n9_adj_8797)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_55_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_35_i5_3_lut (.A(\key_mem[6] [35]), .B(\key_mem[7] [35]), 
         .C(n33952), .Z(n5_adj_8798)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_35_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_55_i8_3_lut (.A(\key_mem[8] [55]), .B(\key_mem[9] [55]), 
         .C(n33952), .Z(n8_adj_8799)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_55_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_55_i5_3_lut (.A(\key_mem[6] [55]), .B(\key_mem[7] [55]), 
         .C(n33952), .Z(n5_adj_8800)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_55_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_55_i4_3_lut (.A(\key_mem[4] [55]), .B(\key_mem[5] [55]), 
         .C(n33952), .Z(n4_adj_8801)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_55_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_35_i4_3_lut (.A(\key_mem[4] [35]), .B(\key_mem[5] [35]), 
         .C(n33952), .Z(n4_adj_8802)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_35_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_35_i2_3_lut (.A(\key_mem[2] [35]), .B(\key_mem[3] [35]), 
         .C(n33952), .Z(n2_adj_8803)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_35_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_55_i2_3_lut (.A(\key_mem[2] [55]), .B(\key_mem[3] [55]), 
         .C(n33952), .Z(n2_adj_8804)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_55_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_35_i1_3_lut (.A(\key_mem[0] [35]), .B(\key_mem[1] [35]), 
         .C(n33952), .Z(n1_adj_8805)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_35_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_55_i1_3_lut (.A(\key_mem[0] [55]), .B(\key_mem[1] [55]), 
         .C(n33952), .Z(n1_adj_8806)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_55_i1_3_lut.init = 16'hcaca;
    LUT4 i15009_2_lut_4_lut (.A(\key_reg[5] [6]), .B(n33655), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[70])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15009_2_lut_4_lut.init = 16'hca00;
    LUT4 round_3__I_0_Mux_54_i11_3_lut (.A(\key_mem[12] [54]), .B(\key_mem[13] [54]), 
         .C(n33952), .Z(n11_adj_64)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_54_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_54_i9_3_lut (.A(\key_mem[10] [54]), .B(\key_mem[11] [54]), 
         .C(n33952), .Z(n9_adj_8808)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_54_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_54_i8_3_lut (.A(\key_mem[8] [54]), .B(\key_mem[9] [54]), 
         .C(n33952), .Z(n8_adj_8809)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_54_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_34_i11_3_lut (.A(\key_mem[12] [34]), .B(\key_mem[13] [34]), 
         .C(n33952), .Z(n11_adj_65)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_34_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_54_i5_3_lut (.A(\key_mem[6] [54]), .B(\key_mem[7] [54]), 
         .C(n33952), .Z(n5_adj_8811)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_54_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_54_i4_3_lut (.A(\key_mem[4] [54]), .B(\key_mem[5] [54]), 
         .C(n33952), .Z(n4_adj_8812)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_54_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_54_i2_3_lut (.A(\key_mem[2] [54]), .B(\key_mem[3] [54]), 
         .C(n33952), .Z(n2_adj_8813)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_54_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_34_i9_3_lut (.A(\key_mem[10] [34]), .B(\key_mem[11] [34]), 
         .C(n33952), .Z(n9_adj_8814)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_34_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_54_i1_3_lut (.A(\key_mem[0] [54]), .B(\key_mem[1] [54]), 
         .C(n33952), .Z(n1_adj_8815)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_54_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_34_i8_3_lut (.A(\key_mem[8] [34]), .B(\key_mem[9] [34]), 
         .C(n33952), .Z(n8_adj_8816)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_34_i8_3_lut.init = 16'hcaca;
    LUT4 i15008_2_lut_4_lut (.A(\key_reg[5] [5]), .B(n33657), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[69])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15008_2_lut_4_lut.init = 16'hca00;
    LUT4 round_3__I_0_Mux_53_i11_3_lut (.A(\key_mem[12] [53]), .B(\key_mem[13] [53]), 
         .C(n33952), .Z(n11_adj_66)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_53_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_34_i5_3_lut (.A(\key_mem[6] [34]), .B(\key_mem[7] [34]), 
         .C(n33952), .Z(n5_adj_8818)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_34_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_53_i9_3_lut (.A(\key_mem[10] [53]), .B(\key_mem[11] [53]), 
         .C(n33952), .Z(n9_adj_8819)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_53_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_53_i8_3_lut (.A(\key_mem[8] [53]), .B(\key_mem[9] [53]), 
         .C(n33952), .Z(n8_adj_8820)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_53_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_34_i4_3_lut (.A(\key_mem[4] [34]), .B(\key_mem[5] [34]), 
         .C(n33952), .Z(n4_adj_8821)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_34_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_34_i2_3_lut (.A(\key_mem[2] [34]), .B(\key_mem[3] [34]), 
         .C(n33952), .Z(n2_adj_8822)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_34_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_53_i5_3_lut (.A(\key_mem[6] [53]), .B(\key_mem[7] [53]), 
         .C(n33952), .Z(n5_adj_8823)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_53_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_34_i1_3_lut (.A(\key_mem[0] [34]), .B(\key_mem[1] [34]), 
         .C(n33952), .Z(n1_adj_8824)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_34_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_53_i4_3_lut (.A(\key_mem[4] [53]), .B(\key_mem[5] [53]), 
         .C(n33952), .Z(n4_adj_8825)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_53_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_53_i2_3_lut (.A(\key_mem[2] [53]), .B(\key_mem[3] [53]), 
         .C(n33952), .Z(n2_adj_8826)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_53_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_53_i1_3_lut (.A(\key_mem[0] [53]), .B(\key_mem[1] [53]), 
         .C(n33952), .Z(n1_adj_8827)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_53_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_33_i11_3_lut (.A(\key_mem[12] [33]), .B(\key_mem[13] [33]), 
         .C(n33952), .Z(n11_adj_67)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_33_i11_3_lut.init = 16'hcaca;
    LUT4 i15007_2_lut_4_lut (.A(\key_reg[5] [4]), .B(n33659), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[68])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15007_2_lut_4_lut.init = 16'hca00;
    LUT4 round_3__I_0_Mux_52_i11_3_lut (.A(\key_mem[12] [52]), .B(\key_mem[13] [52]), 
         .C(n33952), .Z(n11_adj_68)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_52_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_52_i9_3_lut (.A(\key_mem[10] [52]), .B(\key_mem[11] [52]), 
         .C(n33952), .Z(n9_adj_8830)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_52_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_52_i8_3_lut (.A(\key_mem[8] [52]), .B(\key_mem[9] [52]), 
         .C(n33952), .Z(n8_adj_8831)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_52_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_33_i9_3_lut (.A(\key_mem[10] [33]), .B(\key_mem[11] [33]), 
         .C(n33952), .Z(n9_adj_8832)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_33_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_33_i8_3_lut (.A(\key_mem[8] [33]), .B(\key_mem[9] [33]), 
         .C(n33952), .Z(n8_adj_8833)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_33_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_52_i5_3_lut (.A(\key_mem[6] [52]), .B(\key_mem[7] [52]), 
         .C(n33952), .Z(n5_adj_8834)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_52_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_33_i5_3_lut (.A(\key_mem[6] [33]), .B(\key_mem[7] [33]), 
         .C(n33952), .Z(n5_adj_8835)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_33_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_52_i4_3_lut (.A(\key_mem[4] [52]), .B(\key_mem[5] [52]), 
         .C(n33952), .Z(n4_adj_8836)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_52_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_33_i4_3_lut (.A(\key_mem[4] [33]), .B(\key_mem[5] [33]), 
         .C(n33952), .Z(n4_adj_8837)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_33_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_33_i2_3_lut (.A(\key_mem[2] [33]), .B(\key_mem[3] [33]), 
         .C(n33952), .Z(n2_adj_8838)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_33_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_52_i2_3_lut (.A(\key_mem[2] [52]), .B(\key_mem[3] [52]), 
         .C(n33952), .Z(n2_adj_8839)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_52_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_33_i1_3_lut (.A(\key_mem[0] [33]), .B(\key_mem[1] [33]), 
         .C(n33952), .Z(n1_adj_8840)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_33_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_52_i1_3_lut (.A(\key_mem[0] [52]), .B(\key_mem[1] [52]), 
         .C(n33952), .Z(n1_adj_8841)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_52_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_32_i11_3_lut (.A(\key_mem[12] [32]), .B(\key_mem[13] [32]), 
         .C(n33952), .Z(n11_adj_69)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_32_i11_3_lut.init = 16'hcaca;
    LUT4 i15006_2_lut_4_lut (.A(\key_reg[5] [3]), .B(n33661), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[67])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15006_2_lut_4_lut.init = 16'hca00;
    LUT4 round_3__I_0_Mux_32_i9_3_lut (.A(\key_mem[10] [32]), .B(\key_mem[11] [32]), 
         .C(n33952), .Z(n9_adj_8843)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_32_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_51_i11_3_lut (.A(\key_mem[12] [51]), .B(\key_mem[13] [51]), 
         .C(n33952), .Z(n11_adj_70)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_51_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_32_i8_3_lut (.A(\key_mem[8] [32]), .B(\key_mem[9] [32]), 
         .C(n33952), .Z(n8_adj_8845)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_32_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_51_i9_3_lut (.A(\key_mem[10] [51]), .B(\key_mem[11] [51]), 
         .C(n33952), .Z(n9_adj_8846)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_51_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_32_i5_3_lut (.A(\key_mem[6] [32]), .B(\key_mem[7] [32]), 
         .C(n33952), .Z(n5_adj_8847)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_32_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_32_i4_3_lut (.A(\key_mem[4] [32]), .B(\key_mem[5] [32]), 
         .C(n33952), .Z(n4_adj_8848)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_32_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_51_i8_3_lut (.A(\key_mem[8] [51]), .B(\key_mem[9] [51]), 
         .C(n33952), .Z(n8_adj_8849)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_51_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_32_i2_3_lut (.A(\key_mem[2] [32]), .B(\key_mem[3] [32]), 
         .C(n33952), .Z(n2_adj_8850)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_32_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_32_i1_3_lut (.A(\key_mem[0] [32]), .B(\key_mem[1] [32]), 
         .C(n33952), .Z(n1_adj_8851)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_32_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_51_i5_3_lut (.A(\key_mem[6] [51]), .B(\key_mem[7] [51]), 
         .C(n33952), .Z(n5_adj_8852)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_51_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_51_i4_3_lut (.A(\key_mem[4] [51]), .B(\key_mem[5] [51]), 
         .C(n33952), .Z(n4_adj_8853)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_51_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_31_i11_3_lut (.A(\key_mem[12] [31]), .B(\key_mem[13] [31]), 
         .C(n33952), .Z(n11_adj_71)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_31_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_31_i9_3_lut (.A(\key_mem[10] [31]), .B(\key_mem[11] [31]), 
         .C(n33952), .Z(n9_adj_8855)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_31_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_51_i2_3_lut (.A(\key_mem[2] [51]), .B(\key_mem[3] [51]), 
         .C(n33952), .Z(n2_adj_8856)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_51_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_31_i8_3_lut (.A(\key_mem[8] [31]), .B(\key_mem[9] [31]), 
         .C(n33952), .Z(n8_adj_8857)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_31_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_51_i1_3_lut (.A(\key_mem[0] [51]), .B(\key_mem[1] [51]), 
         .C(n33952), .Z(n1_adj_8858)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_51_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_31_i5_3_lut (.A(\key_mem[6] [31]), .B(\key_mem[7] [31]), 
         .C(n33952), .Z(n5_adj_8859)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_31_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_31_i4_3_lut (.A(\key_mem[4] [31]), .B(\key_mem[5] [31]), 
         .C(n33952), .Z(n4_adj_8860)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_31_i4_3_lut.init = 16'hcaca;
    LUT4 i15005_2_lut_4_lut (.A(\key_reg[5] [2]), .B(n33663), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[66])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15005_2_lut_4_lut.init = 16'hca00;
    LUT4 round_3__I_0_Mux_31_i2_3_lut (.A(\key_mem[2] [31]), .B(\key_mem[3] [31]), 
         .C(n33952), .Z(n2_adj_8861)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_31_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_24_i11_3_lut (.A(\key_mem[12] [24]), .B(\key_mem[13] [24]), 
         .C(n33952), .Z(n11_adj_72)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_24_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_31_i1_3_lut (.A(\key_mem[0] [31]), .B(\key_mem[1] [31]), 
         .C(n33952), .Z(n1_adj_8863)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_31_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_24_i9_3_lut (.A(\key_mem[10] [24]), .B(\key_mem[11] [24]), 
         .C(n33952), .Z(n9_adj_8864)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_24_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_30_i11_3_lut (.A(\key_mem[12] [30]), .B(\key_mem[13] [30]), 
         .C(n33952), .Z(n11_adj_73)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_30_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_24_i8_3_lut (.A(\key_mem[8] [24]), .B(\key_mem[9] [24]), 
         .C(n33952), .Z(n8_adj_8866)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_24_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_30_i9_3_lut (.A(\key_mem[10] [30]), .B(\key_mem[11] [30]), 
         .C(n33952), .Z(n9_adj_8867)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_30_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_30_i8_3_lut (.A(\key_mem[8] [30]), .B(\key_mem[9] [30]), 
         .C(n33952), .Z(n8_adj_8868)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_30_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_24_i5_3_lut (.A(\key_mem[6] [24]), .B(\key_mem[7] [24]), 
         .C(n33952), .Z(n5_adj_8869)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_24_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_30_i5_3_lut (.A(\key_mem[6] [30]), .B(\key_mem[7] [30]), 
         .C(n33952), .Z(n5_adj_8870)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_30_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_30_i4_3_lut (.A(\key_mem[4] [30]), .B(\key_mem[5] [30]), 
         .C(n33952), .Z(n4_adj_8871)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_30_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_24_i4_3_lut (.A(\key_mem[4] [24]), .B(\key_mem[5] [24]), 
         .C(n33952), .Z(n4_adj_8872)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_24_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_30_i2_3_lut (.A(\key_mem[2] [30]), .B(\key_mem[3] [30]), 
         .C(n33952), .Z(n2_adj_8873)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_30_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_30_i1_3_lut (.A(\key_mem[0] [30]), .B(\key_mem[1] [30]), 
         .C(n33952), .Z(n1_adj_8874)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_30_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_24_i2_3_lut (.A(\key_mem[2] [24]), .B(\key_mem[3] [24]), 
         .C(n33952), .Z(n2_adj_8875)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_24_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_24_i1_3_lut (.A(\key_mem[0] [24]), .B(\key_mem[1] [24]), 
         .C(n33952), .Z(n1_adj_8876)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_24_i1_3_lut.init = 16'hcaca;
    LUT4 i15004_2_lut_4_lut (.A(\key_reg[5] [1]), .B(n33665), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[65])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15004_2_lut_4_lut.init = 16'hca00;
    LUT4 round_3__I_0_Mux_29_i11_3_lut (.A(\key_mem[12] [29]), .B(\key_mem[13] [29]), 
         .C(n33952), .Z(n11_adj_74)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_29_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_29_i9_3_lut (.A(\key_mem[10] [29]), .B(\key_mem[11] [29]), 
         .C(n33952), .Z(n9_adj_8878)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_29_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_29_i8_3_lut (.A(\key_mem[8] [29]), .B(\key_mem[9] [29]), 
         .C(n33952), .Z(n8_adj_8879)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_29_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_23_i11_3_lut (.A(\key_mem[12] [23]), .B(\key_mem[13] [23]), 
         .C(n33952), .Z(n11_adj_75)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_23_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_29_i5_3_lut (.A(\key_mem[6] [29]), .B(\key_mem[7] [29]), 
         .C(n33952), .Z(n5_adj_8881)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_29_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_29_i4_3_lut (.A(\key_mem[4] [29]), .B(\key_mem[5] [29]), 
         .C(n33952), .Z(n4_adj_8882)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_29_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_23_i9_3_lut (.A(\key_mem[10] [23]), .B(\key_mem[11] [23]), 
         .C(n33952), .Z(n9_adj_8883)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_23_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_29_i2_3_lut (.A(\key_mem[2] [29]), .B(\key_mem[3] [29]), 
         .C(n33952), .Z(n2_adj_8884)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_29_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_29_i1_3_lut (.A(\key_mem[0] [29]), .B(\key_mem[1] [29]), 
         .C(n33952), .Z(n1_adj_8885)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_29_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_23_i8_3_lut (.A(\key_mem[8] [23]), .B(\key_mem[9] [23]), 
         .C(n33952), .Z(n8_adj_8886)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_23_i8_3_lut.init = 16'hcaca;
    LUT4 i15003_2_lut_4_lut (.A(\key_reg[5] [0]), .B(n33666), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[64])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15003_2_lut_4_lut.init = 16'hca00;
    LUT4 round_3__I_0_Mux_28_i11_3_lut (.A(\key_mem[12] [28]), .B(\key_mem[13] [28]), 
         .C(n33952), .Z(n11_adj_76)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_28_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_23_i5_3_lut (.A(\key_mem[6] [23]), .B(\key_mem[7] [23]), 
         .C(n33952), .Z(n5_adj_8888)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_23_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_23_i4_3_lut (.A(\key_mem[4] [23]), .B(\key_mem[5] [23]), 
         .C(n33952), .Z(n4_adj_8889)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_23_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_28_i9_3_lut (.A(\key_mem[10] [28]), .B(\key_mem[11] [28]), 
         .C(n33952), .Z(n9_adj_8890)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_28_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_23_i2_3_lut (.A(\key_mem[2] [23]), .B(\key_mem[3] [23]), 
         .C(n33952), .Z(n2_adj_8891)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_23_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_28_i8_3_lut (.A(\key_mem[8] [28]), .B(\key_mem[9] [28]), 
         .C(n33952), .Z(n8_adj_8892)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_28_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_23_i1_3_lut (.A(\key_mem[0] [23]), .B(\key_mem[1] [23]), 
         .C(n33952), .Z(n1_adj_8893)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_23_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_28_i5_3_lut (.A(\key_mem[6] [28]), .B(\key_mem[7] [28]), 
         .C(n33952), .Z(n5_adj_8894)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_28_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_28_i4_3_lut (.A(\key_mem[4] [28]), .B(\key_mem[5] [28]), 
         .C(n33952), .Z(n4_adj_8895)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_28_i4_3_lut.init = 16'hcaca;
    LUT4 i2_2_lut_rep_254 (.A(prev_key0_reg[95]), .B(n4_adj_8457), .Z(n33558)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i2_2_lut_rep_254.init = 16'h6666;
    LUT4 round_3__I_0_Mux_22_i11_3_lut (.A(\key_mem[12] [22]), .B(\key_mem[13] [22]), 
         .C(n33952), .Z(n11_adj_77)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_22_i11_3_lut.init = 16'hcaca;
    LUT4 i3348_3_lut_4_lut (.A(prev_key1_reg[125]), .B(n33718), .C(n35835), 
         .D(n33528), .Z(n8833)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam i3348_3_lut_4_lut.init = 16'hf606;
    LUT4 round_3__I_0_Mux_28_i2_3_lut (.A(\key_mem[2] [28]), .B(\key_mem[3] [28]), 
         .C(n33952), .Z(n2_adj_8897)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_28_i2_3_lut.init = 16'hcaca;
    L6MUX21 i24994 (.D0(n30151), .D1(n30152), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[43]));
    LUT4 round_3__I_0_Mux_22_i9_3_lut (.A(\key_mem[10] [22]), .B(\key_mem[11] [22]), 
         .C(n33952), .Z(n9_adj_8898)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_22_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_28_i1_3_lut (.A(\key_mem[0] [28]), .B(\key_mem[1] [28]), 
         .C(n33952), .Z(n1_adj_8899)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_28_i1_3_lut.init = 16'hcaca;
    L6MUX21 i25001 (.D0(n30158), .D1(n30159), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[44]));
    LUT4 round_3__I_0_Mux_22_i8_3_lut (.A(\key_mem[8] [22]), .B(\key_mem[9] [22]), 
         .C(n33952), .Z(n8_adj_8900)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_22_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_27_i11_3_lut (.A(\key_mem[12] [27]), .B(\key_mem[13] [27]), 
         .C(n33952), .Z(n11_adj_78)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_27_i11_3_lut.init = 16'hcaca;
    L6MUX21 i25008 (.D0(n30165), .D1(n30166), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[45]));
    LUT4 mux_51_i126_3_lut_4_lut (.A(prev_key1_reg[125]), .B(n33718), .C(n33860), 
         .D(\key_reg[0] [29]), .Z(key_mem_new_127__N_7264[125])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam mux_51_i126_3_lut_4_lut.init = 16'h6f60;
    LUT4 round_3__I_0_Mux_22_i5_3_lut (.A(\key_mem[6] [22]), .B(\key_mem[7] [22]), 
         .C(n33952), .Z(n5_adj_8902)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_22_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_22_i4_3_lut (.A(\key_mem[4] [22]), .B(\key_mem[5] [22]), 
         .C(n33952), .Z(n4_adj_8903)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_22_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_27_i9_3_lut (.A(\key_mem[10] [27]), .B(\key_mem[11] [27]), 
         .C(n33952), .Z(n9_adj_8904)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_27_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_22_i2_3_lut (.A(\key_mem[2] [22]), .B(\key_mem[3] [22]), 
         .C(n33952), .Z(n2_adj_8905)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_22_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_27_i8_3_lut (.A(\key_mem[8] [27]), .B(\key_mem[9] [27]), 
         .C(n33952), .Z(n8_adj_8906)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_27_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_22_i1_3_lut (.A(\key_mem[0] [22]), .B(\key_mem[1] [22]), 
         .C(n33952), .Z(n1_adj_8907)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_22_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_27_i5_3_lut (.A(\key_mem[6] [27]), .B(\key_mem[7] [27]), 
         .C(n33952), .Z(n5_adj_8908)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_27_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_27_i4_3_lut (.A(\key_mem[4] [27]), .B(\key_mem[5] [27]), 
         .C(n33952), .Z(n4_adj_8909)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_27_i4_3_lut.init = 16'hcaca;
    LUT4 mux_85_i96_3_lut_rep_206_4_lut (.A(prev_key0_reg[95]), .B(n4_adj_8457), 
         .C(n33859), .D(\key_reg[5] [31]), .Z(n33510)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam mux_85_i96_3_lut_rep_206_4_lut.init = 16'h6f60;
    L6MUX21 i25015 (.D0(n30172), .D1(n30173), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[46]));
    LUT4 round_3__I_0_Mux_27_i2_3_lut (.A(\key_mem[2] [27]), .B(\key_mem[3] [27]), 
         .C(n33952), .Z(n2_adj_8910)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_27_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_27_i1_3_lut (.A(\key_mem[0] [27]), .B(\key_mem[1] [27]), 
         .C(n33952), .Z(n1_adj_8911)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_27_i1_3_lut.init = 16'hcaca;
    L6MUX21 i25022 (.D0(n30179), .D1(n30180), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[1]));
    LUT4 round_3__I_0_Mux_21_i11_3_lut (.A(\key_mem[12] [21]), .B(\key_mem[13] [21]), 
         .C(n33952), .Z(n11_adj_79)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_21_i11_3_lut.init = 16'hcaca;
    LUT4 i3346_3_lut_4_lut (.A(prev_key1_reg[124]), .B(n33719), .C(n35835), 
         .D(n33529), .Z(n8831)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam i3346_3_lut_4_lut.init = 16'hf606;
    LUT4 round_3__I_0_Mux_25_i11_3_lut (.A(\key_mem[12] [25]), .B(\key_mem[13] [25]), 
         .C(n33952), .Z(n11_adj_80)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_25_i11_3_lut.init = 16'hcaca;
    LUT4 mux_51_i125_3_lut_4_lut (.A(prev_key1_reg[124]), .B(n33719), .C(n33860), 
         .D(\key_reg[0] [28]), .Z(key_mem_new_127__N_7264[124])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam mux_51_i125_3_lut_4_lut.init = 16'h6f60;
    LUT4 round_3__I_0_Mux_21_i9_3_lut (.A(\key_mem[10] [21]), .B(\key_mem[11] [21]), 
         .C(n33952), .Z(n9_adj_8914)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_21_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_25_i9_3_lut (.A(\key_mem[10] [25]), .B(\key_mem[11] [25]), 
         .C(n33952), .Z(n9_adj_8915)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_25_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_21_i8_3_lut (.A(\key_mem[8] [21]), .B(\key_mem[9] [21]), 
         .C(n33952), .Z(n8_adj_8916)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_21_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_25_i8_3_lut (.A(\key_mem[8] [25]), .B(\key_mem[9] [25]), 
         .C(n33952), .Z(n8_adj_8917)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_25_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_25_i5_3_lut (.A(\key_mem[6] [25]), .B(\key_mem[7] [25]), 
         .C(n33952), .Z(n5_adj_8918)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_25_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_25_i4_3_lut (.A(\key_mem[4] [25]), .B(\key_mem[5] [25]), 
         .C(n33952), .Z(n4_adj_8919)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_25_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_21_i5_3_lut (.A(\key_mem[6] [21]), .B(\key_mem[7] [21]), 
         .C(n33952), .Z(n5_adj_8920)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_21_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_127_i11_3_lut (.A(\key_mem[12] [127]), .B(\key_mem[13] [127]), 
         .C(n33952), .Z(n11_adj_81)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_127_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_21_i4_3_lut (.A(\key_mem[4] [21]), .B(\key_mem[5] [21]), 
         .C(n33952), .Z(n4_adj_8922)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_21_i4_3_lut.init = 16'hcaca;
    LUT4 i3344_3_lut_4_lut (.A(prev_key1_reg[123]), .B(n33720), .C(n35835), 
         .D(n33530), .Z(n8829)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam i3344_3_lut_4_lut.init = 16'hf606;
    LUT4 round_3__I_0_Mux_127_i9_3_lut (.A(\key_mem[10] [127]), .B(\key_mem[11] [127]), 
         .C(n33952), .Z(n9_adj_8923)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_127_i9_3_lut.init = 16'hcaca;
    L6MUX21 i25029 (.D0(n30186), .D1(n30187), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[2]));
    LUT4 round_3__I_0_Mux_127_i8_3_lut (.A(\key_mem[8] [127]), .B(\key_mem[9] [127]), 
         .C(n33952), .Z(n8_adj_8924)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_127_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_21_i2_3_lut (.A(\key_mem[2] [21]), .B(\key_mem[3] [21]), 
         .C(n33952), .Z(n2_adj_8925)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_21_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_21_i1_3_lut (.A(\key_mem[0] [21]), .B(\key_mem[1] [21]), 
         .C(n33952), .Z(n1_adj_8926)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_21_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_127_i5_3_lut (.A(\key_mem[6] [127]), .B(\key_mem[7] [127]), 
         .C(n33952), .Z(n5_adj_8927)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_127_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_127_i4_3_lut (.A(\key_mem[4] [127]), .B(\key_mem[5] [127]), 
         .C(n33952), .Z(n4_adj_8928)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_127_i4_3_lut.init = 16'hcaca;
    L6MUX21 i25036 (.D0(n30193), .D1(n30194), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[3]));
    LUT4 round_3__I_0_Mux_20_i11_3_lut (.A(\key_mem[12] [20]), .B(\key_mem[13] [20]), 
         .C(n33952), .Z(n11_adj_82)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_20_i11_3_lut.init = 16'hcaca;
    L6MUX21 i25043 (.D0(n30200), .D1(n30201), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[4]));
    LUT4 mux_51_i124_3_lut_4_lut (.A(prev_key1_reg[123]), .B(n33720), .C(n33860), 
         .D(\key_reg[0] [27]), .Z(key_mem_new_127__N_7264[123])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam mux_51_i124_3_lut_4_lut.init = 16'h6f60;
    LUT4 round_3__I_0_Mux_127_i2_3_lut (.A(\key_mem[2] [127]), .B(\key_mem[3] [127]), 
         .C(n33952), .Z(n2_adj_8930)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_127_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_127_i1_3_lut (.A(\key_mem[0] [127]), .B(\key_mem[1] [127]), 
         .C(n33952), .Z(n1_adj_8931)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_127_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_20_i9_3_lut (.A(\key_mem[10] [20]), .B(\key_mem[11] [20]), 
         .C(n33952), .Z(n9_adj_8932)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_20_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_20_i8_3_lut (.A(\key_mem[8] [20]), .B(\key_mem[9] [20]), 
         .C(n33952), .Z(n8_adj_8933)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_20_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_20_i5_3_lut (.A(\key_mem[6] [20]), .B(\key_mem[7] [20]), 
         .C(n33952), .Z(n5_adj_8934)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_20_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_126_i11_3_lut (.A(\key_mem[12] [126]), .B(\key_mem[13] [126]), 
         .C(n33952), .Z(n11_adj_83)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_126_i11_3_lut.init = 16'hcaca;
    LUT4 i3342_3_lut_4_lut (.A(prev_key1_reg[122]), .B(n33721), .C(n35835), 
         .D(n33531), .Z(n8827)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam i3342_3_lut_4_lut.init = 16'hf606;
    LUT4 round_3__I_0_Mux_20_i4_3_lut (.A(\key_mem[4] [20]), .B(\key_mem[5] [20]), 
         .C(n33952), .Z(n4_adj_8936)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_20_i4_3_lut.init = 16'hcaca;
    L6MUX21 i25050 (.D0(n30207), .D1(n30208), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[5]));
    LUT4 round_3__I_0_Mux_20_i2_3_lut (.A(\key_mem[2] [20]), .B(\key_mem[3] [20]), 
         .C(n33952), .Z(n2_adj_8937)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_20_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_20_i1_3_lut (.A(\key_mem[0] [20]), .B(\key_mem[1] [20]), 
         .C(n33952), .Z(n1_adj_8938)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_20_i1_3_lut.init = 16'hcaca;
    LUT4 i2_2_lut_rep_257 (.A(prev_key0_reg[94]), .B(n4_adj_8455), .Z(n33561)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i2_2_lut_rep_257.init = 16'h6666;
    LUT4 round_3__I_0_Mux_50_i11_3_lut (.A(\key_mem[12] [50]), .B(\key_mem[13] [50]), 
         .C(n33952), .Z(n11_adj_84)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_50_i11_3_lut.init = 16'hcaca;
    LUT4 mux_51_i123_3_lut_4_lut (.A(prev_key1_reg[122]), .B(n33721), .C(n33860), 
         .D(\key_reg[0] [26]), .Z(key_mem_new_127__N_7264[122])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam mux_51_i123_3_lut_4_lut.init = 16'h6f60;
    L6MUX21 i25057 (.D0(n30214), .D1(n30215), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[6]));
    LUT4 round_3__I_0_Mux_50_i9_3_lut (.A(\key_mem[10] [50]), .B(\key_mem[11] [50]), 
         .C(n33952), .Z(n9_adj_8940)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_50_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_126_i9_3_lut (.A(\key_mem[10] [126]), .B(\key_mem[11] [126]), 
         .C(n33952), .Z(n9_adj_8941)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_126_i9_3_lut.init = 16'hcaca;
    L6MUX21 i25064 (.D0(n30221), .D1(n30222), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[26]));
    L6MUX21 i25071 (.D0(n30228), .D1(n30229), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[7]));
    LUT4 round_3__I_0_Mux_50_i8_3_lut (.A(\key_mem[8] [50]), .B(\key_mem[9] [50]), 
         .C(n33952), .Z(n8_adj_8942)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_50_i8_3_lut.init = 16'hcaca;
    L6MUX21 i25078 (.D0(n30235), .D1(n30236), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[8]));
    L6MUX21 i25085 (.D0(n30242), .D1(n30243), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[0]));
    LUT4 round_3__I_0_Mux_50_i5_3_lut (.A(\key_mem[6] [50]), .B(\key_mem[7] [50]), 
         .C(n33952), .Z(n5_adj_8943)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_50_i5_3_lut.init = 16'hcaca;
    L6MUX21 i25092 (.D0(n30249), .D1(n30250), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[9]));
    L6MUX21 i25099 (.D0(n30256), .D1(n30257), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[10]));
    LUT4 round_3__I_0_Mux_50_i4_3_lut (.A(\key_mem[4] [50]), .B(\key_mem[5] [50]), 
         .C(n33952), .Z(n4_adj_8944)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_50_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_50_i2_3_lut (.A(\key_mem[2] [50]), .B(\key_mem[3] [50]), 
         .C(n33952), .Z(n2_adj_8945)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_50_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_50_i1_3_lut (.A(\key_mem[0] [50]), .B(\key_mem[1] [50]), 
         .C(n33952), .Z(n1_adj_8946)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_50_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_126_i8_3_lut (.A(\key_mem[8] [126]), .B(\key_mem[9] [126]), 
         .C(n33952), .Z(n8_adj_8947)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_126_i8_3_lut.init = 16'hcaca;
    L6MUX21 i25106 (.D0(n30263), .D1(n30264), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[11]));
    LUT4 round_3__I_0_Mux_19_i11_3_lut (.A(\key_mem[12] [19]), .B(\key_mem[13] [19]), 
         .C(n33952), .Z(n11_adj_85)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_19_i11_3_lut.init = 16'hcaca;
    L6MUX21 i25113 (.D0(n30270), .D1(n30271), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[12]));
    L6MUX21 i25120 (.D0(n30277), .D1(n30278), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[13]));
    LUT4 i3338_3_lut_4_lut (.A(prev_key1_reg[120]), .B(n33723), .C(n35835), 
         .D(n33533), .Z(n8823)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam i3338_3_lut_4_lut.init = 16'hf606;
    LUT4 round_3__I_0_Mux_19_i9_3_lut (.A(\key_mem[10] [19]), .B(\key_mem[11] [19]), 
         .C(n33952), .Z(n9_adj_8949)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_19_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_19_i8_3_lut (.A(\key_mem[8] [19]), .B(\key_mem[9] [19]), 
         .C(n33952), .Z(n8_adj_8950)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_19_i8_3_lut.init = 16'hcaca;
    L6MUX21 i25127 (.D0(n30284), .D1(n30285), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[14]));
    LUT4 round_3__I_0_Mux_19_i5_3_lut (.A(\key_mem[6] [19]), .B(\key_mem[7] [19]), 
         .C(n33952), .Z(n5_adj_8951)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_19_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_126_i5_3_lut (.A(\key_mem[6] [126]), .B(\key_mem[7] [126]), 
         .C(n33952), .Z(n5_adj_8952)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_126_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_126_i4_3_lut (.A(\key_mem[4] [126]), .B(\key_mem[5] [126]), 
         .C(n33952), .Z(n4_adj_8953)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_126_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_19_i4_3_lut (.A(\key_mem[4] [19]), .B(\key_mem[5] [19]), 
         .C(n33952), .Z(n4_adj_8954)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_19_i4_3_lut.init = 16'hcaca;
    L6MUX21 i25134 (.D0(n30291), .D1(n30292), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[15]));
    L6MUX21 i25141 (.D0(n30298), .D1(n30299), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[16]));
    L6MUX21 i25148 (.D0(n30305), .D1(n30306), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[47]));
    L6MUX21 i25155 (.D0(n30312), .D1(n30313), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[48]));
    L6MUX21 i25162 (.D0(n30319), .D1(n30320), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[49]));
    L6MUX21 i25169 (.D0(n30326), .D1(n30327), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[17]));
    LUT4 round_3__I_0_Mux_126_i2_3_lut (.A(\key_mem[2] [126]), .B(\key_mem[3] [126]), 
         .C(n33952), .Z(n2_adj_8955)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_126_i2_3_lut.init = 16'hcaca;
    PFUMX i25682 (.BLUT(n4_adj_8956), .ALUT(n5_adj_8957), .C0(\muxed_round_nr[1] ), 
          .Z(n30841));
    L6MUX21 i25176 (.D0(n30333), .D1(n30334), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[18]));
    LUT4 round_3__I_0_Mux_126_i1_3_lut (.A(\key_mem[0] [126]), .B(\key_mem[1] [126]), 
         .C(n33952), .Z(n1_adj_8958)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_126_i1_3_lut.init = 16'hcaca;
    LUT4 mux_85_i95_3_lut_rep_207_4_lut (.A(prev_key0_reg[94]), .B(n4_adj_8455), 
         .C(n33859), .D(\key_reg[5] [30]), .Z(n33511)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam mux_85_i95_3_lut_rep_207_4_lut.init = 16'h6f60;
    LUT4 round_3__I_0_Mux_19_i2_3_lut (.A(\key_mem[2] [19]), .B(\key_mem[3] [19]), 
         .C(n33952), .Z(n2_adj_8959)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_19_i2_3_lut.init = 16'hcaca;
    L6MUX21 i25183 (.D0(n30340), .D1(n30341), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[19]));
    LUT4 round_3__I_0_Mux_19_i1_3_lut (.A(\key_mem[0] [19]), .B(\key_mem[1] [19]), 
         .C(n33952), .Z(n1_adj_8960)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_19_i1_3_lut.init = 16'hcaca;
    LUT4 i2_2_lut_rep_258 (.A(prev_key0_reg[93]), .B(n4_adj_8451), .Z(n33562)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i2_2_lut_rep_258.init = 16'h6666;
    L6MUX21 i25190 (.D0(n30347), .D1(n30348), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[50]));
    LUT4 round_3__I_0_Mux_18_i11_3_lut (.A(\key_mem[12] [18]), .B(\key_mem[13] [18]), 
         .C(n33952), .Z(n11_adj_86)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_18_i11_3_lut.init = 16'hcaca;
    LUT4 mux_51_i121_3_lut_4_lut (.A(prev_key1_reg[120]), .B(n33723), .C(n33860), 
         .D(\key_reg[0] [24]), .Z(key_mem_new_127__N_7264[120])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam mux_51_i121_3_lut_4_lut.init = 16'h6f60;
    LUT4 round_3__I_0_Mux_18_i9_3_lut (.A(\key_mem[10] [18]), .B(\key_mem[11] [18]), 
         .C(n33952), .Z(n9_adj_8962)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_18_i9_3_lut.init = 16'hcaca;
    L6MUX21 i25197 (.D0(n30354), .D1(n30355), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[20]));
    L6MUX21 i25204 (.D0(n30361), .D1(n30362), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[21]));
    L6MUX21 i25211 (.D0(n30368), .D1(n30369), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[22]));
    L6MUX21 i25218 (.D0(n30375), .D1(n30376), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[23]));
    LUT4 round_3__I_0_Mux_18_i8_3_lut (.A(\key_mem[8] [18]), .B(\key_mem[9] [18]), 
         .C(n33952), .Z(n8_adj_8963)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_18_i8_3_lut.init = 16'hcaca;
    L6MUX21 i25225 (.D0(n30382), .D1(n30383), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[24]));
    LUT4 round_3__I_0_Mux_18_i5_3_lut (.A(\key_mem[6] [18]), .B(\key_mem[7] [18]), 
         .C(n33952), .Z(n5_adj_8964)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_18_i5_3_lut.init = 16'hcaca;
    L6MUX21 i25232 (.D0(n30389), .D1(n30390), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[51]));
    L6MUX21 i25239 (.D0(n30396), .D1(n30397), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[52]));
    LUT4 round_3__I_0_Mux_18_i4_3_lut (.A(\key_mem[4] [18]), .B(\key_mem[5] [18]), 
         .C(n33952), .Z(n4_adj_8965)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_18_i4_3_lut.init = 16'hcaca;
    L6MUX21 i25246 (.D0(n30403), .D1(n30404), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[53]));
    LUT4 round_3__I_0_Mux_18_i2_3_lut (.A(\key_mem[2] [18]), .B(\key_mem[3] [18]), 
         .C(n33952), .Z(n2_adj_8966)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_18_i2_3_lut.init = 16'hcaca;
    L6MUX21 i25253 (.D0(n30410), .D1(n30411), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[54]));
    L6MUX21 i25260 (.D0(n30417), .D1(n30418), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[55]));
    LUT4 round_3__I_0_Mux_18_i1_3_lut (.A(\key_mem[0] [18]), .B(\key_mem[1] [18]), 
         .C(n33952), .Z(n1_adj_8967)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_18_i1_3_lut.init = 16'hcaca;
    L6MUX21 i25267 (.D0(n30424), .D1(n30425), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[56]));
    L6MUX21 i25274 (.D0(n30431), .D1(n30432), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[57]));
    L6MUX21 i25281 (.D0(n30438), .D1(n30439), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[58]));
    L6MUX21 i25288 (.D0(n30445), .D1(n30446), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[59]));
    L6MUX21 i25295 (.D0(n30452), .D1(n30453), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[60]));
    LUT4 round_3__I_0_Mux_125_i11_3_lut (.A(\key_mem[12] [125]), .B(\key_mem[13] [125]), 
         .C(n33952), .Z(n11_adj_87)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_125_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_17_i11_3_lut (.A(\key_mem[12] [17]), .B(\key_mem[13] [17]), 
         .C(n33952), .Z(n11_adj_88)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_17_i11_3_lut.init = 16'hcaca;
    L6MUX21 i25302 (.D0(n30459), .D1(n30460), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[61]));
    L6MUX21 i25309 (.D0(n30466), .D1(n30467), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[62]));
    LUT4 round_3__I_0_Mux_17_i9_3_lut (.A(\key_mem[10] [17]), .B(\key_mem[11] [17]), 
         .C(n33952), .Z(n9_adj_8970)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_17_i9_3_lut.init = 16'hcaca;
    L6MUX21 i25316 (.D0(n30473), .D1(n30474), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[63]));
    L6MUX21 i25323 (.D0(n30480), .D1(n30481), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[64]));
    LUT4 round_3__I_0_Mux_17_i8_3_lut (.A(\key_mem[8] [17]), .B(\key_mem[9] [17]), 
         .C(n33952), .Z(n8_adj_8971)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_17_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_17_i5_3_lut (.A(\key_mem[6] [17]), .B(\key_mem[7] [17]), 
         .C(n33952), .Z(n5_adj_8972)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_17_i5_3_lut.init = 16'hcaca;
    L6MUX21 i25330 (.D0(n30487), .D1(n30488), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[65]));
    L6MUX21 i25337 (.D0(n30494), .D1(n30495), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[66]));
    L6MUX21 i25344 (.D0(n30501), .D1(n30502), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[67]));
    LUT4 round_3__I_0_Mux_17_i4_3_lut (.A(\key_mem[4] [17]), .B(\key_mem[5] [17]), 
         .C(n33952), .Z(n4_adj_8973)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_17_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_17_i2_3_lut (.A(\key_mem[2] [17]), .B(\key_mem[3] [17]), 
         .C(n33952), .Z(n2_adj_8974)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_17_i2_3_lut.init = 16'hcaca;
    LUT4 i15058_2_lut_4_lut (.A(\key_reg[4] [23]), .B(n4_adj_8421), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[119])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15058_2_lut_4_lut.init = 16'hca00;
    LUT4 round_3__I_0_Mux_17_i1_3_lut (.A(\key_mem[0] [17]), .B(\key_mem[1] [17]), 
         .C(n33952), .Z(n1_adj_8975)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_17_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_125_i9_3_lut (.A(\key_mem[10] [125]), .B(\key_mem[11] [125]), 
         .C(n33952), .Z(n9_adj_8976)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_125_i9_3_lut.init = 16'hcaca;
    LUT4 mux_85_i94_3_lut_rep_208_4_lut (.A(prev_key0_reg[93]), .B(n4_adj_8451), 
         .C(n33859), .D(\key_reg[5] [29]), .Z(n33512)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam mux_85_i94_3_lut_rep_208_4_lut.init = 16'h6f60;
    LUT4 round_3__I_0_Mux_125_i8_3_lut (.A(\key_mem[8] [125]), .B(\key_mem[9] [125]), 
         .C(n33952), .Z(n8_adj_8977)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_125_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_49_i11_3_lut (.A(\key_mem[12] [49]), .B(\key_mem[13] [49]), 
         .C(n33952), .Z(n11_adj_89)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_49_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_49_i9_3_lut (.A(\key_mem[10] [49]), .B(\key_mem[11] [49]), 
         .C(n33952), .Z(n9_adj_8979)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_49_i9_3_lut.init = 16'hcaca;
    LUT4 i11158_4_lut (.A(\key_reg[7] [23]), .B(n33621), .C(n33859), .D(n4_adj_8980), 
         .Z(n16742)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i11158_4_lut.init = 16'h3aca;
    LUT4 round_3__I_0_Mux_49_i8_3_lut (.A(\key_mem[8] [49]), .B(\key_mem[9] [49]), 
         .C(n33952), .Z(n8_adj_8981)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_49_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_49_i5_3_lut (.A(\key_mem[6] [49]), .B(\key_mem[7] [49]), 
         .C(n33952), .Z(n5_adj_8982)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_49_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_49_i4_3_lut (.A(\key_mem[4] [49]), .B(\key_mem[5] [49]), 
         .C(n33952), .Z(n4_adj_8983)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_49_i4_3_lut.init = 16'hcaca;
    LUT4 i11097_4_lut (.A(\key_reg[7] [22]), .B(n33623), .C(n33859), .D(n4_adj_8984), 
         .Z(n16682)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i11097_4_lut.init = 16'h3aca;
    LUT4 round_3__I_0_Mux_49_i2_3_lut (.A(\key_mem[2] [49]), .B(\key_mem[3] [49]), 
         .C(n33952), .Z(n2_adj_8985)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_49_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_125_i5_3_lut (.A(\key_mem[6] [125]), .B(\key_mem[7] [125]), 
         .C(n33952), .Z(n5_adj_8986)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_125_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_49_i1_3_lut (.A(\key_mem[0] [49]), .B(\key_mem[1] [49]), 
         .C(n33952), .Z(n1_adj_8987)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_49_i1_3_lut.init = 16'hcaca;
    LUT4 i11036_4_lut (.A(\key_reg[7] [21]), .B(n33625), .C(n33859), .D(n4_adj_8988), 
         .Z(n16622)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i11036_4_lut.init = 16'h3aca;
    LUT4 round_3__I_0_Mux_48_i11_3_lut (.A(\key_mem[12] [48]), .B(\key_mem[13] [48]), 
         .C(n33952), .Z(n11_adj_90)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_48_i11_3_lut.init = 16'hcaca;
    LUT4 i10975_4_lut (.A(\key_reg[7] [20]), .B(n33627), .C(n33859), .D(n4_adj_8990), 
         .Z(n16562)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i10975_4_lut.init = 16'h3aca;
    LUT4 i15057_2_lut_4_lut (.A(\key_reg[4] [22]), .B(n4_adj_8417), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[118])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15057_2_lut_4_lut.init = 16'hca00;
    LUT4 round_3__I_0_Mux_125_i4_3_lut (.A(\key_mem[4] [125]), .B(\key_mem[5] [125]), 
         .C(n33952), .Z(n4_adj_8991)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_125_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_48_i9_3_lut (.A(\key_mem[10] [48]), .B(\key_mem[11] [48]), 
         .C(n33952), .Z(n9_adj_8992)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_48_i9_3_lut.init = 16'hcaca;
    LUT4 i10914_4_lut (.A(\key_reg[7] [19]), .B(n33629), .C(n33859), .D(n4_adj_8993), 
         .Z(n16502)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i10914_4_lut.init = 16'h3aca;
    LUT4 round_3__I_0_Mux_48_i8_3_lut (.A(\key_mem[8] [48]), .B(\key_mem[9] [48]), 
         .C(n33952), .Z(n8_adj_8994)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_48_i8_3_lut.init = 16'hcaca;
    LUT4 i10853_4_lut (.A(\key_reg[7] [18]), .B(n33631), .C(n33859), .D(n4_adj_8995), 
         .Z(n16442)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i10853_4_lut.init = 16'h3aca;
    LUT4 round_3__I_0_Mux_48_i5_3_lut (.A(\key_mem[6] [48]), .B(\key_mem[7] [48]), 
         .C(n33952), .Z(n5_adj_8996)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_48_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_48_i4_3_lut (.A(\key_mem[4] [48]), .B(\key_mem[5] [48]), 
         .C(n33952), .Z(n4_adj_8997)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_48_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_48_i2_3_lut (.A(\key_mem[2] [48]), .B(\key_mem[3] [48]), 
         .C(n33952), .Z(n2_adj_8998)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_48_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_48_i1_3_lut (.A(\key_mem[0] [48]), .B(\key_mem[1] [48]), 
         .C(n33952), .Z(n1_adj_8999)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_48_i1_3_lut.init = 16'hcaca;
    LUT4 i10792_4_lut (.A(\key_reg[7] [17]), .B(n33633), .C(n33859), .D(n4_adj_9000), 
         .Z(n16382)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i10792_4_lut.init = 16'h3aca;
    LUT4 i10731_4_lut (.A(\key_reg[7] [16]), .B(n33635), .C(n33859), .D(n4_adj_9001), 
         .Z(n16322)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i10731_4_lut.init = 16'h3aca;
    LUT4 round_3__I_0_Mux_125_i2_3_lut (.A(\key_mem[2] [125]), .B(\key_mem[3] [125]), 
         .C(n33952), .Z(n2_adj_9002)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_125_i2_3_lut.init = 16'hcaca;
    LUT4 i6_2_lut_3_lut_adj_617 (.A(prev_key1_reg[61]), .B(n33615), .C(keymem_sboxw[29]), 
         .Z(n17097)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;
    defparam i6_2_lut_3_lut_adj_617.init = 16'h9696;
    LUT4 i10670_4_lut (.A(\key_reg[7] [15]), .B(n33637), .C(n33859), .D(n4_adj_9003), 
         .Z(n16262)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i10670_4_lut.init = 16'h3aca;
    LUT4 round_3__I_0_Mux_47_i11_3_lut (.A(\key_mem[12] [47]), .B(\key_mem[13] [47]), 
         .C(n33952), .Z(n11_adj_91)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_47_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_125_i1_3_lut (.A(\key_mem[0] [125]), .B(\key_mem[1] [125]), 
         .C(n33952), .Z(n1_adj_9005)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_125_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_47_i9_3_lut (.A(\key_mem[10] [47]), .B(\key_mem[11] [47]), 
         .C(n33952), .Z(n9_adj_9006)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_47_i9_3_lut.init = 16'hcaca;
    LUT4 i10609_4_lut (.A(\key_reg[7] [14]), .B(n33639), .C(n33859), .D(n4_adj_9007), 
         .Z(n16202)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i10609_4_lut.init = 16'h3aca;
    LUT4 round_3__I_0_Mux_47_i8_3_lut (.A(\key_mem[8] [47]), .B(\key_mem[9] [47]), 
         .C(n33952), .Z(n8_adj_9008)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_47_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_47_i5_3_lut (.A(\key_mem[6] [47]), .B(\key_mem[7] [47]), 
         .C(n33952), .Z(n5_adj_9009)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_47_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_47_i4_3_lut (.A(\key_mem[4] [47]), .B(\key_mem[5] [47]), 
         .C(n33952), .Z(n4_adj_9010)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_47_i4_3_lut.init = 16'hcaca;
    LUT4 i10548_4_lut (.A(\key_reg[7] [13]), .B(n33641), .C(n33859), .D(n4_adj_9011), 
         .Z(n16142)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i10548_4_lut.init = 16'h3aca;
    LUT4 round_3__I_0_Mux_47_i2_3_lut (.A(\key_mem[2] [47]), .B(\key_mem[3] [47]), 
         .C(n33952), .Z(n2_adj_9012)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_47_i2_3_lut.init = 16'hcaca;
    LUT4 i10487_4_lut (.A(\key_reg[7] [12]), .B(n33643), .C(n33859), .D(n4_adj_9013), 
         .Z(n16082)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i10487_4_lut.init = 16'h3aca;
    LUT4 round_3__I_0_Mux_47_i1_3_lut (.A(\key_mem[0] [47]), .B(\key_mem[1] [47]), 
         .C(n33952), .Z(n1_adj_9014)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_47_i1_3_lut.init = 16'hcaca;
    LUT4 i6_2_lut_3_lut_adj_618 (.A(prev_key1_reg[60]), .B(n33616), .C(keymem_sboxw[28]), 
         .Z(n17037)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;
    defparam i6_2_lut_3_lut_adj_618.init = 16'h9696;
    LUT4 i10426_4_lut (.A(\key_reg[7] [11]), .B(n33645), .C(n33859), .D(n4_adj_9015), 
         .Z(n16022)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i10426_4_lut.init = 16'h3aca;
    LUT4 round_3__I_0_Mux_16_i11_3_lut (.A(\key_mem[12] [16]), .B(\key_mem[13] [16]), 
         .C(n33952), .Z(n11_adj_92)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_16_i11_3_lut.init = 16'hcaca;
    LUT4 i15056_2_lut_4_lut (.A(\key_reg[4] [21]), .B(n4_adj_8410), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[117])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15056_2_lut_4_lut.init = 16'hca00;
    LUT4 round_3__I_0_Mux_16_i9_3_lut (.A(\key_mem[10] [16]), .B(\key_mem[11] [16]), 
         .C(n33952), .Z(n9_adj_9017)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_16_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_16_i8_3_lut (.A(\key_mem[8] [16]), .B(\key_mem[9] [16]), 
         .C(n33952), .Z(n8_adj_9018)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_16_i8_3_lut.init = 16'hcaca;
    LUT4 i10365_4_lut (.A(\key_reg[7] [10]), .B(n33647), .C(n33859), .D(n4_adj_9019), 
         .Z(n15962)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i10365_4_lut.init = 16'h3aca;
    L6MUX21 i25351 (.D0(n30508), .D1(n30509), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[68]));
    L6MUX21 i25358 (.D0(n30515), .D1(n30516), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[69]));
    LUT4 round_3__I_0_Mux_124_i11_3_lut (.A(\key_mem[12] [124]), .B(\key_mem[13] [124]), 
         .C(n33952), .Z(n11_adj_93)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_124_i11_3_lut.init = 16'hcaca;
    LUT4 i10304_4_lut (.A(\key_reg[7] [9]), .B(n33649), .C(n33859), .D(n4_adj_9021), 
         .Z(n15902)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i10304_4_lut.init = 16'h3aca;
    LUT4 round_3__I_0_Mux_16_i5_3_lut (.A(\key_mem[6] [16]), .B(\key_mem[7] [16]), 
         .C(n33952), .Z(n5_adj_9022)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_16_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_16_i4_3_lut (.A(\key_mem[4] [16]), .B(\key_mem[5] [16]), 
         .C(n33952), .Z(n4_adj_9023)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_16_i4_3_lut.init = 16'hcaca;
    LUT4 i10243_4_lut (.A(\key_reg[7] [8]), .B(n33651), .C(n33859), .D(n4_adj_9024), 
         .Z(n15842)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i10243_4_lut.init = 16'h3aca;
    LUT4 round_3__I_0_Mux_16_i2_3_lut (.A(\key_mem[2] [16]), .B(\key_mem[3] [16]), 
         .C(n33952), .Z(n2_adj_9025)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_16_i2_3_lut.init = 16'hcaca;
    L6MUX21 i25365 (.D0(n30522), .D1(n30523), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[70]));
    L6MUX21 i25372 (.D0(n30529), .D1(n30530), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[71]));
    L6MUX21 i25379 (.D0(n30536), .D1(n30537), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[72]));
    L6MUX21 i25386 (.D0(n30543), .D1(n30544), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[73]));
    L6MUX21 i25393 (.D0(n30550), .D1(n30551), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[74]));
    L6MUX21 i25400 (.D0(n30557), .D1(n30558), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[75]));
    L6MUX21 i25407 (.D0(n30564), .D1(n30565), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[76]));
    L6MUX21 i25414 (.D0(n30571), .D1(n30572), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[77]));
    L6MUX21 i25421 (.D0(n30578), .D1(n30579), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[78]));
    L6MUX21 i25428 (.D0(n30585), .D1(n30586), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[79]));
    L6MUX21 i25435 (.D0(n30592), .D1(n30593), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[80]));
    LUT4 round_3__I_0_Mux_16_i1_3_lut (.A(\key_mem[0] [16]), .B(\key_mem[1] [16]), 
         .C(n33952), .Z(n1_adj_9026)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_16_i1_3_lut.init = 16'hcaca;
    LUT4 i10182_4_lut (.A(\key_reg[7] [7]), .B(n33653), .C(n33859), .D(n4_adj_9027), 
         .Z(n15782)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i10182_4_lut.init = 16'h3aca;
    L6MUX21 i25442 (.D0(n30599), .D1(n30600), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[81]));
    L6MUX21 i25449 (.D0(n30606), .D1(n30607), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[82]));
    LUT4 i2_2_lut_rep_261 (.A(prev_key0_reg[92]), .B(n4_adj_8449), .Z(n33565)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i2_2_lut_rep_261.init = 16'h6666;
    L6MUX21 i25456 (.D0(n30613), .D1(n30614), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[83]));
    LUT4 round_3__I_0_Mux_15_i11_3_lut (.A(\key_mem[12] [15]), .B(\key_mem[13] [15]), 
         .C(n33952), .Z(n11_adj_94)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_15_i11_3_lut.init = 16'hcaca;
    L6MUX21 i25463 (.D0(n30620), .D1(n30621), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[84]));
    LUT4 i10121_4_lut (.A(\key_reg[7] [6]), .B(n33655), .C(n33859), .D(n4_adj_9029), 
         .Z(n15722)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i10121_4_lut.init = 16'h3aca;
    LUT4 i15055_2_lut_4_lut (.A(\key_reg[4] [20]), .B(n4_adj_8403), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[116])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15055_2_lut_4_lut.init = 16'hca00;
    L6MUX21 i25470 (.D0(n30627), .D1(n30628), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[85]));
    LUT4 round_3__I_0_Mux_15_i9_3_lut (.A(\key_mem[10] [15]), .B(\key_mem[11] [15]), 
         .C(n33952), .Z(n9_adj_9030)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_15_i9_3_lut.init = 16'hcaca;
    L6MUX21 i25477 (.D0(n30634), .D1(n30635), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[86]));
    LUT4 round_3__I_0_Mux_15_i8_3_lut (.A(\key_mem[8] [15]), .B(\key_mem[9] [15]), 
         .C(n33952), .Z(n8_adj_9031)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_15_i8_3_lut.init = 16'hcaca;
    L6MUX21 i25484 (.D0(n30641), .D1(n30642), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[87]));
    L6MUX21 i25491 (.D0(n30648), .D1(n30649), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[88]));
    L6MUX21 i25498 (.D0(n30655), .D1(n30656), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[89]));
    L6MUX21 i25505 (.D0(n30662), .D1(n30663), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[90]));
    L6MUX21 i25512 (.D0(n30669), .D1(n30670), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[91]));
    L6MUX21 i25519 (.D0(n30676), .D1(n30677), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[92]));
    L6MUX21 i25526 (.D0(n30683), .D1(n30684), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[93]));
    L6MUX21 i25533 (.D0(n30690), .D1(n30691), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[94]));
    L6MUX21 i25540 (.D0(n30697), .D1(n30698), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[95]));
    L6MUX21 i25547 (.D0(n30704), .D1(n30705), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[96]));
    L6MUX21 i25554 (.D0(n30711), .D1(n30712), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[97]));
    LUT4 i10060_4_lut (.A(\key_reg[7] [5]), .B(n33657), .C(n33859), .D(n4_adj_9032), 
         .Z(n15662)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i10060_4_lut.init = 16'h3aca;
    L6MUX21 i25561 (.D0(n30718), .D1(n30719), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[98]));
    L6MUX21 i25568 (.D0(n30725), .D1(n30726), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[99]));
    L6MUX21 i25575 (.D0(n30732), .D1(n30733), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[100]));
    LUT4 round_3__I_0_Mux_15_i5_3_lut (.A(\key_mem[6] [15]), .B(\key_mem[7] [15]), 
         .C(n33952), .Z(n5_adj_9033)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_15_i5_3_lut.init = 16'hcaca;
    L6MUX21 i25582 (.D0(n30739), .D1(n30740), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[101]));
    L6MUX21 i25589 (.D0(n30746), .D1(n30747), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[102]));
    L6MUX21 i25596 (.D0(n30753), .D1(n30754), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[103]));
    L6MUX21 i25603 (.D0(n30760), .D1(n30761), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[104]));
    L6MUX21 i25610 (.D0(n30767), .D1(n30768), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[105]));
    L6MUX21 i25617 (.D0(n30774), .D1(n30775), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[106]));
    L6MUX21 i25624 (.D0(n30781), .D1(n30782), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[107]));
    L6MUX21 i25631 (.D0(n30788), .D1(n30789), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[108]));
    L6MUX21 i25638 (.D0(n30795), .D1(n30796), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[109]));
    L6MUX21 i25645 (.D0(n30802), .D1(n30803), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[110]));
    L6MUX21 i25652 (.D0(n30809), .D1(n30810), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[111]));
    LUT4 i9999_4_lut (.A(\key_reg[7] [4]), .B(n33659), .C(n33859), .D(n4_adj_9034), 
         .Z(n15602)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i9999_4_lut.init = 16'h3aca;
    L6MUX21 i25659 (.D0(n30816), .D1(n30817), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[112]));
    L6MUX21 i25666 (.D0(n30823), .D1(n30824), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[113]));
    L6MUX21 i25673 (.D0(n30830), .D1(n30831), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[114]));
    LUT4 round_3__I_0_Mux_15_i4_3_lut (.A(\key_mem[4] [15]), .B(\key_mem[5] [15]), 
         .C(n33952), .Z(n4_adj_9035)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_15_i4_3_lut.init = 16'hcaca;
    L6MUX21 i25680 (.D0(n30837), .D1(n30838), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[115]));
    LUT4 round_3__I_0_Mux_124_i9_3_lut (.A(\key_mem[10] [124]), .B(\key_mem[11] [124]), 
         .C(n33952), .Z(n9_adj_9036)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_124_i9_3_lut.init = 16'hcaca;
    L6MUX21 i25687 (.D0(n30844), .D1(n30845), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[116]));
    LUT4 round_3__I_0_Mux_124_i8_3_lut (.A(\key_mem[8] [124]), .B(\key_mem[9] [124]), 
         .C(n33952), .Z(n8_adj_9037)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_124_i8_3_lut.init = 16'hcaca;
    L6MUX21 i25694 (.D0(n30851), .D1(n30852), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[117]));
    L6MUX21 i25701 (.D0(n30858), .D1(n30859), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[118]));
    L6MUX21 i25708 (.D0(n30865), .D1(n30866), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[119]));
    LUT4 round_3__I_0_Mux_15_i2_3_lut (.A(\key_mem[2] [15]), .B(\key_mem[3] [15]), 
         .C(n33952), .Z(n2_adj_9038)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_15_i2_3_lut.init = 16'hcaca;
    L6MUX21 i25715 (.D0(n30872), .D1(n30873), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[120]));
    L6MUX21 i25722 (.D0(n30879), .D1(n30880), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[121]));
    LUT4 round_3__I_0_Mux_15_i1_3_lut (.A(\key_mem[0] [15]), .B(\key_mem[1] [15]), 
         .C(n33952), .Z(n1_adj_9039)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_15_i1_3_lut.init = 16'hcaca;
    L6MUX21 i25729 (.D0(n30886), .D1(n30887), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[122]));
    L6MUX21 i25736 (.D0(n30893), .D1(n30894), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[123]));
    L6MUX21 i25743 (.D0(n30900), .D1(n30901), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[124]));
    L6MUX21 i25750 (.D0(n30907), .D1(n30908), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[125]));
    L6MUX21 i25757 (.D0(n30914), .D1(n30915), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[126]));
    L6MUX21 i25764 (.D0(n30921), .D1(n30922), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[127]));
    LUT4 i9938_4_lut (.A(\key_reg[7] [3]), .B(n33661), .C(n33859), .D(n4_adj_9040), 
         .Z(n15542)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i9938_4_lut.init = 16'h3aca;
    L6MUX21 i25867 (.D0(n31024), .D1(n31025), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[25]));
    L6MUX21 i25874 (.D0(n31031), .D1(n31032), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[27]));
    L6MUX21 i25881 (.D0(n31038), .D1(n31039), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[28]));
    L6MUX21 i25888 (.D0(n31045), .D1(n31046), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[29]));
    L6MUX21 i25895 (.D0(n31052), .D1(n31053), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[30]));
    L6MUX21 i25902 (.D0(n31059), .D1(n31060), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[31]));
    L6MUX21 i25909 (.D0(n31066), .D1(n31067), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[32]));
    L6MUX21 i25916 (.D0(n31073), .D1(n31074), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[33]));
    L6MUX21 i25923 (.D0(n31080), .D1(n31081), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[34]));
    L6MUX21 i25930 (.D0(n31087), .D1(n31088), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[35]));
    L6MUX21 i25937 (.D0(n31094), .D1(n31095), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[36]));
    L6MUX21 i25944 (.D0(n31101), .D1(n31102), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[37]));
    L6MUX21 i25951 (.D0(n31108), .D1(n31109), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[38]));
    L6MUX21 i25958 (.D0(n31115), .D1(n31116), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[39]));
    L6MUX21 i25965 (.D0(n31122), .D1(n31123), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[40]));
    L6MUX21 i25972 (.D0(n31129), .D1(n31130), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[41]));
    L6MUX21 i25979 (.D0(n31136), .D1(n31137), .SD(\muxed_round_nr[3] ), 
            .Z(round_key[42]));
    LUT4 round_3__I_0_Mux_14_i11_3_lut (.A(\key_mem[12] [14]), .B(\key_mem[13] [14]), 
         .C(n33952), .Z(n11_adj_95)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_14_i11_3_lut.init = 16'hcaca;
    L6MUX21 i24992 (.D0(n30147), .D1(n30148), .SD(\muxed_round_nr[2] ), 
            .Z(n30151));
    LUT4 i9877_4_lut (.A(\key_reg[7] [2]), .B(n33663), .C(n33859), .D(n4_adj_9042), 
         .Z(n15482)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i9877_4_lut.init = 16'h3aca;
    L6MUX21 i24993 (.D0(n30149), .D1(n33343), .SD(\muxed_round_nr[2] ), 
            .Z(n30152));
    LUT4 round_3__I_0_Mux_14_i9_3_lut (.A(\key_mem[10] [14]), .B(\key_mem[11] [14]), 
         .C(n33952), .Z(n9_adj_9043)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_14_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_124_i5_3_lut (.A(\key_mem[6] [124]), .B(\key_mem[7] [124]), 
         .C(n33952), .Z(n5_adj_9044)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_124_i5_3_lut.init = 16'hcaca;
    L6MUX21 i24999 (.D0(n30154), .D1(n30155), .SD(\muxed_round_nr[2] ), 
            .Z(n30158));
    L6MUX21 i25000 (.D0(n30156), .D1(n33344), .SD(\muxed_round_nr[2] ), 
            .Z(n30159));
    L6MUX21 i25006 (.D0(n30161), .D1(n30162), .SD(\muxed_round_nr[2] ), 
            .Z(n30165));
    L6MUX21 i25007 (.D0(n30163), .D1(n33345), .SD(\muxed_round_nr[2] ), 
            .Z(n30166));
    LUT4 round_3__I_0_Mux_124_i4_3_lut (.A(\key_mem[4] [124]), .B(\key_mem[5] [124]), 
         .C(n33952), .Z(n4_adj_9045)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_124_i4_3_lut.init = 16'hcaca;
    L6MUX21 i25013 (.D0(n30168), .D1(n30169), .SD(\muxed_round_nr[2] ), 
            .Z(n30172));
    L6MUX21 i25014 (.D0(n30170), .D1(n33346), .SD(\muxed_round_nr[2] ), 
            .Z(n30173));
    LUT4 i9816_4_lut (.A(\key_reg[7] [1]), .B(n33665), .C(n33859), .D(n4_adj_9046), 
         .Z(n15422)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i9816_4_lut.init = 16'h3aca;
    L6MUX21 i25020 (.D0(n30175), .D1(n30176), .SD(\muxed_round_nr[2] ), 
            .Z(n30179));
    L6MUX21 i25021 (.D0(n30177), .D1(n33347), .SD(\muxed_round_nr[2] ), 
            .Z(n30180));
    L6MUX21 i25027 (.D0(n30182), .D1(n30183), .SD(\muxed_round_nr[2] ), 
            .Z(n30186));
    L6MUX21 i25028 (.D0(n30184), .D1(n33348), .SD(\muxed_round_nr[2] ), 
            .Z(n30187));
    L6MUX21 i25034 (.D0(n30189), .D1(n30190), .SD(\muxed_round_nr[2] ), 
            .Z(n30193));
    L6MUX21 i25035 (.D0(n30191), .D1(n33349), .SD(\muxed_round_nr[2] ), 
            .Z(n30194));
    L6MUX21 i25041 (.D0(n30196), .D1(n30197), .SD(\muxed_round_nr[2] ), 
            .Z(n30200));
    L6MUX21 i25042 (.D0(n30198), .D1(n33351), .SD(\muxed_round_nr[2] ), 
            .Z(n30201));
    L6MUX21 i25048 (.D0(n30203), .D1(n30204), .SD(\muxed_round_nr[2] ), 
            .Z(n30207));
    L6MUX21 i25049 (.D0(n30205), .D1(n33352), .SD(\muxed_round_nr[2] ), 
            .Z(n30208));
    L6MUX21 i25055 (.D0(n30210), .D1(n30211), .SD(\muxed_round_nr[2] ), 
            .Z(n30214));
    L6MUX21 i25056 (.D0(n30212), .D1(n33353), .SD(\muxed_round_nr[2] ), 
            .Z(n30215));
    L6MUX21 i25062 (.D0(n30217), .D1(n30218), .SD(\muxed_round_nr[2] ), 
            .Z(n30221));
    L6MUX21 i25063 (.D0(n30219), .D1(n33354), .SD(\muxed_round_nr[2] ), 
            .Z(n30222));
    L6MUX21 i25069 (.D0(n30224), .D1(n30225), .SD(\muxed_round_nr[2] ), 
            .Z(n30228));
    L6MUX21 i25070 (.D0(n30226), .D1(n33356), .SD(\muxed_round_nr[2] ), 
            .Z(n30229));
    L6MUX21 i25076 (.D0(n30231), .D1(n30232), .SD(\muxed_round_nr[2] ), 
            .Z(n30235));
    L6MUX21 i25077 (.D0(n30233), .D1(n33357), .SD(\muxed_round_nr[2] ), 
            .Z(n30236));
    L6MUX21 i25083 (.D0(n30238), .D1(n30239), .SD(\muxed_round_nr[2] ), 
            .Z(n30242));
    LUT4 round_3__I_0_Mux_14_i8_3_lut (.A(\key_mem[8] [14]), .B(\key_mem[9] [14]), 
         .C(n33952), .Z(n8_adj_9047)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_14_i8_3_lut.init = 16'hcaca;
    L6MUX21 i25084 (.D0(n30240), .D1(n33358), .SD(\muxed_round_nr[2] ), 
            .Z(n30243));
    L6MUX21 i25090 (.D0(n30245), .D1(n30246), .SD(\muxed_round_nr[2] ), 
            .Z(n30249));
    LUT4 i9701_4_lut (.A(\key_reg[7] [0]), .B(n33666), .C(n33859), .D(n4_adj_9048), 
         .Z(n15309)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i9701_4_lut.init = 16'h3aca;
    L6MUX21 i25091 (.D0(n30247), .D1(n33359), .SD(\muxed_round_nr[2] ), 
            .Z(n30250));
    LUT4 round_3__I_0_Mux_14_i5_3_lut (.A(\key_mem[6] [14]), .B(\key_mem[7] [14]), 
         .C(n33952), .Z(n5_adj_9049)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_14_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_14_i4_3_lut (.A(\key_mem[4] [14]), .B(\key_mem[5] [14]), 
         .C(n33952), .Z(n4_adj_9050)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_14_i4_3_lut.init = 16'hcaca;
    L6MUX21 i25097 (.D0(n30252), .D1(n30253), .SD(\muxed_round_nr[2] ), 
            .Z(n30256));
    LUT4 i11646_4_lut (.A(\key_reg[7] [31]), .B(n33558), .C(n33859), .D(n4_adj_9051), 
         .Z(n17222)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i11646_4_lut.init = 16'h3aca;
    LUT4 round_3__I_0_Mux_14_i2_3_lut (.A(\key_mem[2] [14]), .B(\key_mem[3] [14]), 
         .C(n33952), .Z(n2_adj_9052)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_14_i2_3_lut.init = 16'hcaca;
    L6MUX21 i25098 (.D0(n30254), .D1(n33360), .SD(\muxed_round_nr[2] ), 
            .Z(n30257));
    LUT4 round_3__I_0_Mux_14_i1_3_lut (.A(\key_mem[0] [14]), .B(\key_mem[1] [14]), 
         .C(n33952), .Z(n1_adj_9053)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_14_i1_3_lut.init = 16'hcaca;
    L6MUX21 i25104 (.D0(n30259), .D1(n30260), .SD(\muxed_round_nr[2] ), 
            .Z(n30263));
    L6MUX21 i25105 (.D0(n30261), .D1(n33362), .SD(\muxed_round_nr[2] ), 
            .Z(n30264));
    L6MUX21 i25111 (.D0(n30266), .D1(n30267), .SD(\muxed_round_nr[2] ), 
            .Z(n30270));
    L6MUX21 i25112 (.D0(n30268), .D1(n33363), .SD(\muxed_round_nr[2] ), 
            .Z(n30271));
    L6MUX21 i25118 (.D0(n30273), .D1(n30274), .SD(\muxed_round_nr[2] ), 
            .Z(n30277));
    L6MUX21 i25119 (.D0(n30275), .D1(n33364), .SD(\muxed_round_nr[2] ), 
            .Z(n30278));
    LUT4 mux_85_i93_3_lut_rep_209_4_lut (.A(prev_key0_reg[92]), .B(n4_adj_8449), 
         .C(n33859), .D(\key_reg[5] [28]), .Z(n33513)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam mux_85_i93_3_lut_rep_209_4_lut.init = 16'h6f60;
    L6MUX21 i25125 (.D0(n30280), .D1(n30281), .SD(\muxed_round_nr[2] ), 
            .Z(n30284));
    L6MUX21 i25126 (.D0(n30282), .D1(n33365), .SD(\muxed_round_nr[2] ), 
            .Z(n30285));
    L6MUX21 i25132 (.D0(n30287), .D1(n30288), .SD(\muxed_round_nr[2] ), 
            .Z(n30291));
    LUT4 i11585_4_lut (.A(\key_reg[7] [30]), .B(n33561), .C(n33859), .D(n4_adj_9054), 
         .Z(n17162)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i11585_4_lut.init = 16'h3aca;
    LUT4 i11524_4_lut (.A(\key_reg[7] [29]), .B(n33562), .C(n33859), .D(n4_adj_9055), 
         .Z(n17102)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i11524_4_lut.init = 16'h3aca;
    LUT4 round_3__I_0_Mux_13_i11_3_lut (.A(\key_mem[12] [13]), .B(\key_mem[13] [13]), 
         .C(n33952), .Z(n11_adj_96)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_13_i11_3_lut.init = 16'hcaca;
    LUT4 i15054_2_lut_4_lut (.A(\key_reg[4] [19]), .B(n4_adj_8400), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[115])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15054_2_lut_4_lut.init = 16'hca00;
    LUT4 round_3__I_0_Mux_13_i9_3_lut (.A(\key_mem[10] [13]), .B(\key_mem[11] [13]), 
         .C(n33952), .Z(n9_adj_9057)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_13_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_13_i8_3_lut (.A(\key_mem[8] [13]), .B(\key_mem[9] [13]), 
         .C(n33952), .Z(n8_adj_9058)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_13_i8_3_lut.init = 16'hcaca;
    LUT4 i11463_4_lut (.A(\key_reg[7] [28]), .B(n33565), .C(n33859), .D(n4_adj_9059), 
         .Z(n17042)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i11463_4_lut.init = 16'h3aca;
    LUT4 round_3__I_0_Mux_13_i5_3_lut (.A(\key_mem[6] [13]), .B(\key_mem[7] [13]), 
         .C(n33952), .Z(n5_adj_9060)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_13_i5_3_lut.init = 16'hcaca;
    LUT4 i11402_4_lut (.A(\key_reg[7] [27]), .B(n33567), .C(n33859), .D(n4_adj_9061), 
         .Z(n16982)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i11402_4_lut.init = 16'h3aca;
    L6MUX21 i25133 (.D0(n30289), .D1(n33366), .SD(\muxed_round_nr[2] ), 
            .Z(n30292));
    L6MUX21 i25139 (.D0(n30294), .D1(n30295), .SD(\muxed_round_nr[2] ), 
            .Z(n30298));
    L6MUX21 i25140 (.D0(n30296), .D1(n33368), .SD(\muxed_round_nr[2] ), 
            .Z(n30299));
    L6MUX21 i25146 (.D0(n30301), .D1(n30302), .SD(\muxed_round_nr[2] ), 
            .Z(n30305));
    L6MUX21 i25147 (.D0(n30303), .D1(n33369), .SD(\muxed_round_nr[2] ), 
            .Z(n30306));
    L6MUX21 i25153 (.D0(n30308), .D1(n30309), .SD(\muxed_round_nr[2] ), 
            .Z(n30312));
    L6MUX21 i25154 (.D0(n30310), .D1(n33370), .SD(\muxed_round_nr[2] ), 
            .Z(n30313));
    LUT4 round_3__I_0_Mux_13_i4_3_lut (.A(\key_mem[4] [13]), .B(\key_mem[5] [13]), 
         .C(n33952), .Z(n4_adj_9062)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_13_i4_3_lut.init = 16'hcaca;
    L6MUX21 i25160 (.D0(n30315), .D1(n30316), .SD(\muxed_round_nr[2] ), 
            .Z(n30319));
    L6MUX21 i25161 (.D0(n30317), .D1(n33371), .SD(\muxed_round_nr[2] ), 
            .Z(n30320));
    L6MUX21 i25167 (.D0(n30322), .D1(n30323), .SD(\muxed_round_nr[2] ), 
            .Z(n30326));
    LUT4 round_3__I_0_Mux_13_i2_3_lut (.A(\key_mem[2] [13]), .B(\key_mem[3] [13]), 
         .C(n33952), .Z(n2_adj_9063)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_13_i2_3_lut.init = 16'hcaca;
    LUT4 i11341_4_lut (.A(\key_reg[7] [26]), .B(n33568), .C(n33859), .D(n4_adj_9064), 
         .Z(n16922)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i11341_4_lut.init = 16'h3aca;
    LUT4 round_3__I_0_Mux_13_i1_3_lut (.A(\key_mem[0] [13]), .B(\key_mem[1] [13]), 
         .C(n33952), .Z(n1_adj_9065)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_13_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_12_i11_3_lut (.A(\key_mem[12] [12]), .B(\key_mem[13] [12]), 
         .C(n33952), .Z(n11_adj_97)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_12_i11_3_lut.init = 16'hcaca;
    LUT4 i11280_4_lut (.A(\key_reg[7] [25]), .B(n33571), .C(n33859), .D(n4_adj_9067), 
         .Z(n16862)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i11280_4_lut.init = 16'h3aca;
    LUT4 round_3__I_0_Mux_12_i9_3_lut (.A(\key_mem[10] [12]), .B(\key_mem[11] [12]), 
         .C(n33952), .Z(n9_adj_9068)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_12_i9_3_lut.init = 16'hcaca;
    L6MUX21 i25168 (.D0(n30324), .D1(n33372), .SD(\muxed_round_nr[2] ), 
            .Z(n30327));
    L6MUX21 i25174 (.D0(n30329), .D1(n30330), .SD(\muxed_round_nr[2] ), 
            .Z(n30333));
    L6MUX21 i25175 (.D0(n30331), .D1(n33373), .SD(\muxed_round_nr[2] ), 
            .Z(n30334));
    L6MUX21 i25181 (.D0(n30336), .D1(n30337), .SD(\muxed_round_nr[2] ), 
            .Z(n30340));
    L6MUX21 i25182 (.D0(n30338), .D1(n33375), .SD(\muxed_round_nr[2] ), 
            .Z(n30341));
    LUT4 round_3__I_0_Mux_12_i8_3_lut (.A(\key_mem[8] [12]), .B(\key_mem[9] [12]), 
         .C(n33952), .Z(n8_adj_9069)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_12_i8_3_lut.init = 16'hcaca;
    L6MUX21 i25188 (.D0(n30343), .D1(n30344), .SD(\muxed_round_nr[2] ), 
            .Z(n30347));
    L6MUX21 i25189 (.D0(n30345), .D1(n33376), .SD(\muxed_round_nr[2] ), 
            .Z(n30348));
    LUT4 i1_3_lut_4_lut (.A(n33860), .B(\key_reg[3] [0]), .C(n15311), 
         .D(n35839), .Z(key_mem_new[0])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_3_lut_4_lut.init = 16'hf400;
    L6MUX21 i25195 (.D0(n30350), .D1(n30351), .SD(\muxed_round_nr[2] ), 
            .Z(n30354));
    LUT4 i1_3_lut_4_lut_adj_619 (.A(n33860), .B(\key_reg[3] [0]), .C(n15311), 
         .D(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[0])) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_3_lut_4_lut_adj_619.init = 16'hf0f4;
    L6MUX21 i25196 (.D0(n30352), .D1(n33378), .SD(\muxed_round_nr[2] ), 
            .Z(n30355));
    L6MUX21 i25202 (.D0(n30357), .D1(n30358), .SD(\muxed_round_nr[2] ), 
            .Z(n30361));
    LUT4 round_3__I_0_Mux_12_i5_3_lut (.A(\key_mem[6] [12]), .B(\key_mem[7] [12]), 
         .C(n33952), .Z(n5_adj_9070)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_12_i5_3_lut.init = 16'hcaca;
    L6MUX21 i25203 (.D0(n30359), .D1(n33381), .SD(\muxed_round_nr[2] ), 
            .Z(n30362));
    LUT4 round_3__I_0_Mux_12_i4_3_lut (.A(\key_mem[4] [12]), .B(\key_mem[5] [12]), 
         .C(n33952), .Z(n4_adj_9071)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_12_i4_3_lut.init = 16'hcaca;
    L6MUX21 i25209 (.D0(n30364), .D1(n30365), .SD(\muxed_round_nr[2] ), 
            .Z(n30368));
    LUT4 round_3__I_0_Mux_12_i2_3_lut (.A(\key_mem[2] [12]), .B(\key_mem[3] [12]), 
         .C(n33952), .Z(n2_adj_9072)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_12_i2_3_lut.init = 16'hcaca;
    L6MUX21 i25210 (.D0(n30366), .D1(n33383), .SD(\muxed_round_nr[2] ), 
            .Z(n30369));
    LUT4 round_3__I_0_Mux_12_i1_3_lut (.A(\key_mem[0] [12]), .B(\key_mem[1] [12]), 
         .C(n33952), .Z(n1_adj_9073)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_12_i1_3_lut.init = 16'hcaca;
    L6MUX21 i25216 (.D0(n30371), .D1(n30372), .SD(\muxed_round_nr[2] ), 
            .Z(n30375));
    L6MUX21 i25217 (.D0(n30373), .D1(n33385), .SD(\muxed_round_nr[2] ), 
            .Z(n30376));
    L6MUX21 i25223 (.D0(n30378), .D1(n30379), .SD(\muxed_round_nr[2] ), 
            .Z(n30382));
    L6MUX21 i25224 (.D0(n30380), .D1(n33388), .SD(\muxed_round_nr[2] ), 
            .Z(n30383));
    L6MUX21 i25230 (.D0(n30385), .D1(n30386), .SD(\muxed_round_nr[2] ), 
            .Z(n30389));
    L6MUX21 i25231 (.D0(n30387), .D1(n33390), .SD(\muxed_round_nr[2] ), 
            .Z(n30390));
    L6MUX21 i25237 (.D0(n30392), .D1(n30393), .SD(\muxed_round_nr[2] ), 
            .Z(n30396));
    LUT4 i6_2_lut_3_lut_adj_620 (.A(prev_key1_reg[59]), .B(n33617), .C(keymem_sboxw[27]), 
         .Z(n16977)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;
    defparam i6_2_lut_3_lut_adj_620.init = 16'h9696;
    LUT4 round_3__I_0_Mux_11_i11_3_lut (.A(\key_mem[12] [11]), .B(\key_mem[13] [11]), 
         .C(n33952), .Z(n11_adj_98)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_11_i11_3_lut.init = 16'hcaca;
    LUT4 i15053_2_lut_4_lut (.A(\key_reg[4] [18]), .B(n4_adj_8395), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[114])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15053_2_lut_4_lut.init = 16'hca00;
    LUT4 round_3__I_0_Mux_11_i9_3_lut (.A(\key_mem[10] [11]), .B(\key_mem[11] [11]), 
         .C(n33952), .Z(n9_adj_9075)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_11_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_11_i8_3_lut (.A(\key_mem[8] [11]), .B(\key_mem[9] [11]), 
         .C(n33952), .Z(n8_adj_9076)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_11_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_11_i5_3_lut (.A(\key_mem[6] [11]), .B(\key_mem[7] [11]), 
         .C(n33952), .Z(n5_adj_9077)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_11_i5_3_lut.init = 16'hcaca;
    LUT4 i15098_3_lut_4_lut (.A(n33860), .B(\key_reg[2] [31]), .C(n17229), 
         .D(n35839), .Z(key_mem_new[63])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i15098_3_lut_4_lut.init = 16'hf400;
    LUT4 round_3__I_0_Mux_124_i2_3_lut (.A(\key_mem[2] [124]), .B(\key_mem[3] [124]), 
         .C(n33952), .Z(n2_adj_9078)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_124_i2_3_lut.init = 16'hcaca;
    LUT4 i15097_3_lut_4_lut (.A(n33860), .B(\key_reg[2] [30]), .C(n17169), 
         .D(n35839), .Z(key_mem_new[62])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i15097_3_lut_4_lut.init = 16'hf400;
    LUT4 round_3__I_0_Mux_11_i4_3_lut (.A(\key_mem[4] [11]), .B(\key_mem[5] [11]), 
         .C(n33952), .Z(n4_adj_9079)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_11_i4_3_lut.init = 16'hcaca;
    LUT4 i15096_3_lut_4_lut (.A(n33860), .B(\key_reg[2] [29]), .C(n17109), 
         .D(n35839), .Z(key_mem_new[61])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i15096_3_lut_4_lut.init = 16'hf400;
    LUT4 i15095_3_lut_4_lut (.A(n33860), .B(\key_reg[2] [28]), .C(n17049), 
         .D(n35839), .Z(key_mem_new[60])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i15095_3_lut_4_lut.init = 16'hf400;
    LUT4 round_3__I_0_Mux_124_i1_3_lut (.A(\key_mem[0] [124]), .B(\key_mem[1] [124]), 
         .C(n33952), .Z(n1_adj_9080)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_124_i1_3_lut.init = 16'hcaca;
    LUT4 i15094_3_lut_4_lut (.A(n33860), .B(\key_reg[2] [27]), .C(n16989), 
         .D(n35839), .Z(key_mem_new[59])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i15094_3_lut_4_lut.init = 16'hf400;
    LUT4 i15093_3_lut_4_lut (.A(n33860), .B(\key_reg[2] [26]), .C(n16929), 
         .D(n35839), .Z(key_mem_new[58])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i15093_3_lut_4_lut.init = 16'hf400;
    LUT4 round_3__I_0_Mux_11_i2_3_lut (.A(\key_mem[2] [11]), .B(\key_mem[3] [11]), 
         .C(n33952), .Z(n2_adj_9081)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_11_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_11_i1_3_lut (.A(\key_mem[0] [11]), .B(\key_mem[1] [11]), 
         .C(n33952), .Z(n1_adj_9082)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_11_i1_3_lut.init = 16'hcaca;
    LUT4 i15092_3_lut_4_lut (.A(n33860), .B(\key_reg[2] [25]), .C(n16869), 
         .D(n35839), .Z(key_mem_new[57])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i15092_3_lut_4_lut.init = 16'hf400;
    LUT4 i15091_3_lut_4_lut (.A(n33860), .B(\key_reg[2] [24]), .C(n16809), 
         .D(n35839), .Z(key_mem_new[56])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i15091_3_lut_4_lut.init = 16'hf400;
    LUT4 i2_2_lut_rep_263 (.A(prev_key0_reg[91]), .B(n4_adj_8444), .Z(n33567)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i2_2_lut_rep_263.init = 16'h6666;
    LUT4 round_3__I_0_Mux_10_i11_3_lut (.A(\key_mem[12] [10]), .B(\key_mem[13] [10]), 
         .C(n33952), .Z(n11_adj_99)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_10_i11_3_lut.init = 16'hcaca;
    LUT4 i15090_3_lut_4_lut (.A(n33860), .B(\key_reg[2] [23]), .C(n16749), 
         .D(n35839), .Z(key_mem_new[55])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i15090_3_lut_4_lut.init = 16'hf400;
    LUT4 i15089_3_lut_4_lut (.A(n33860), .B(\key_reg[2] [22]), .C(n16689), 
         .D(n35839), .Z(key_mem_new[54])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i15089_3_lut_4_lut.init = 16'hf400;
    LUT4 i15088_3_lut_4_lut (.A(n33860), .B(\key_reg[2] [21]), .C(n16629), 
         .D(n35839), .Z(key_mem_new[53])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i15088_3_lut_4_lut.init = 16'hf400;
    LUT4 i11219_4_lut (.A(\key_reg[7] [24]), .B(n33573), .C(n33859), .D(n4_adj_9084), 
         .Z(n16802)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(81[17:29])
    defparam i11219_4_lut.init = 16'h3aca;
    LUT4 i15087_3_lut_4_lut (.A(n33860), .B(\key_reg[2] [20]), .C(n16569), 
         .D(n35839), .Z(key_mem_new[52])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i15087_3_lut_4_lut.init = 16'hf400;
    LUT4 i15086_3_lut_4_lut (.A(n33860), .B(\key_reg[2] [19]), .C(n16509), 
         .D(n35839), .Z(key_mem_new[51])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i15086_3_lut_4_lut.init = 16'hf400;
    LUT4 i15085_3_lut_4_lut (.A(n33860), .B(\key_reg[2] [18]), .C(n16449), 
         .D(n35839), .Z(key_mem_new[50])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i15085_3_lut_4_lut.init = 16'hf400;
    LUT4 round_3__I_0_Mux_10_i9_3_lut (.A(\key_mem[10] [10]), .B(\key_mem[11] [10]), 
         .C(n33952), .Z(n9_adj_9085)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_10_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_10_i8_3_lut (.A(\key_mem[8] [10]), .B(\key_mem[9] [10]), 
         .C(n33952), .Z(n8_adj_9086)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_10_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_10_i5_3_lut (.A(\key_mem[6] [10]), .B(\key_mem[7] [10]), 
         .C(n33952), .Z(n5_adj_9087)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_10_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_10_i4_3_lut (.A(\key_mem[4] [10]), .B(\key_mem[5] [10]), 
         .C(n33952), .Z(n4_adj_9088)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_10_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_10_i2_3_lut (.A(\key_mem[2] [10]), .B(\key_mem[3] [10]), 
         .C(n33952), .Z(n2_adj_9089)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_10_i2_3_lut.init = 16'hcaca;
    LUT4 i15084_3_lut_4_lut (.A(n33860), .B(\key_reg[2] [17]), .C(n16389), 
         .D(n35839), .Z(key_mem_new[49])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i15084_3_lut_4_lut.init = 16'hf400;
    LUT4 i15083_3_lut_4_lut (.A(n33860), .B(\key_reg[2] [16]), .C(n16329), 
         .D(n35839), .Z(key_mem_new[48])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i15083_3_lut_4_lut.init = 16'hf400;
    LUT4 i15082_3_lut_4_lut (.A(n33860), .B(\key_reg[2] [15]), .C(n16269), 
         .D(n35839), .Z(key_mem_new[47])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i15082_3_lut_4_lut.init = 16'hf400;
    LUT4 round_3__I_0_Mux_123_i11_3_lut (.A(\key_mem[12] [123]), .B(\key_mem[13] [123]), 
         .C(n33952), .Z(n11_adj_100)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_123_i11_3_lut.init = 16'hcaca;
    LUT4 i15081_3_lut_4_lut (.A(n33860), .B(\key_reg[2] [14]), .C(n16209), 
         .D(n35839), .Z(key_mem_new[46])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i15081_3_lut_4_lut.init = 16'hf400;
    LUT4 i15052_2_lut_4_lut (.A(\key_reg[4] [17]), .B(n4_adj_8390), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[113])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15052_2_lut_4_lut.init = 16'hca00;
    L6MUX21 i25238 (.D0(n30394), .D1(n33392), .SD(\muxed_round_nr[2] ), 
            .Z(n30397));
    LUT4 i15080_3_lut_4_lut (.A(n33860), .B(\key_reg[2] [13]), .C(n16149), 
         .D(n35839), .Z(key_mem_new[45])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i15080_3_lut_4_lut.init = 16'hf400;
    LUT4 round_3__I_0_Mux_10_i1_3_lut (.A(\key_mem[0] [10]), .B(\key_mem[1] [10]), 
         .C(n33952), .Z(n1_adj_9091)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_10_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_123_i9_3_lut (.A(\key_mem[10] [123]), .B(\key_mem[11] [123]), 
         .C(n33952), .Z(n9_adj_9092)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_123_i9_3_lut.init = 16'hcaca;
    LUT4 i15079_3_lut_4_lut (.A(n33860), .B(\key_reg[2] [12]), .C(n16089), 
         .D(n35839), .Z(key_mem_new[44])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i15079_3_lut_4_lut.init = 16'hf400;
    LUT4 round_3__I_0_Mux_123_i8_3_lut (.A(\key_mem[8] [123]), .B(\key_mem[9] [123]), 
         .C(n33952), .Z(n8_adj_9093)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_123_i8_3_lut.init = 16'hcaca;
    LUT4 mux_85_i92_3_lut_rep_210_4_lut (.A(prev_key0_reg[91]), .B(n4_adj_8444), 
         .C(n33859), .D(\key_reg[5] [27]), .Z(n33514)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam mux_85_i92_3_lut_rep_210_4_lut.init = 16'h6f60;
    LUT4 round_3__I_0_Mux_9_i11_3_lut (.A(\key_mem[12] [9]), .B(\key_mem[13] [9]), 
         .C(n33952), .Z(n11_adj_101)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_9_i11_3_lut.init = 16'hcaca;
    LUT4 i15078_3_lut_4_lut (.A(n33860), .B(\key_reg[2] [11]), .C(n16029), 
         .D(n35839), .Z(key_mem_new[43])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i15078_3_lut_4_lut.init = 16'hf400;
    LUT4 i15077_3_lut_4_lut (.A(n33860), .B(\key_reg[2] [10]), .C(n15969), 
         .D(n35839), .Z(key_mem_new[42])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i15077_3_lut_4_lut.init = 16'hf400;
    LUT4 i15076_3_lut_4_lut (.A(n33860), .B(\key_reg[2] [9]), .C(n15909), 
         .D(n35839), .Z(key_mem_new[41])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i15076_3_lut_4_lut.init = 16'hf400;
    LUT4 round_3__I_0_Mux_9_i9_3_lut (.A(\key_mem[10] [9]), .B(\key_mem[11] [9]), 
         .C(n33952), .Z(n9_adj_9095)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_9_i9_3_lut.init = 16'hcaca;
    LUT4 i15075_3_lut_4_lut (.A(n33860), .B(\key_reg[2] [8]), .C(n15849), 
         .D(n35839), .Z(key_mem_new[40])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i15075_3_lut_4_lut.init = 16'hf400;
    LUT4 i15074_3_lut_4_lut (.A(n33860), .B(\key_reg[2] [7]), .C(n15789), 
         .D(n35839), .Z(key_mem_new[39])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i15074_3_lut_4_lut.init = 16'hf400;
    LUT4 i15073_3_lut_4_lut (.A(n33860), .B(\key_reg[2] [6]), .C(n15729), 
         .D(n35839), .Z(key_mem_new[38])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i15073_3_lut_4_lut.init = 16'hf400;
    LUT4 round_3__I_0_Mux_9_i8_3_lut (.A(\key_mem[8] [9]), .B(\key_mem[9] [9]), 
         .C(n33952), .Z(n8_adj_9096)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_9_i8_3_lut.init = 16'hcaca;
    LUT4 i15072_3_lut_4_lut (.A(n33860), .B(\key_reg[2] [5]), .C(n15669), 
         .D(n35839), .Z(key_mem_new[37])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i15072_3_lut_4_lut.init = 16'hf400;
    LUT4 i15071_3_lut_4_lut (.A(n33860), .B(\key_reg[2] [4]), .C(n15609), 
         .D(n35839), .Z(key_mem_new[36])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i15071_3_lut_4_lut.init = 16'hf400;
    LUT4 round_3__I_0_Mux_9_i5_3_lut (.A(\key_mem[6] [9]), .B(\key_mem[7] [9]), 
         .C(n33952), .Z(n5_adj_9097)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_9_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_9_i4_3_lut (.A(\key_mem[4] [9]), .B(\key_mem[5] [9]), 
         .C(n33952), .Z(n4_adj_9098)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_9_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_9_i2_3_lut (.A(\key_mem[2] [9]), .B(\key_mem[3] [9]), 
         .C(n33952), .Z(n2_adj_9099)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_9_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_9_i1_3_lut (.A(\key_mem[0] [9]), .B(\key_mem[1] [9]), 
         .C(n33952), .Z(n1_adj_9100)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_9_i1_3_lut.init = 16'hcaca;
    LUT4 i15070_3_lut_4_lut (.A(n33860), .B(\key_reg[2] [3]), .C(n15549), 
         .D(n35839), .Z(key_mem_new[35])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i15070_3_lut_4_lut.init = 16'hf400;
    LUT4 i15069_3_lut_4_lut (.A(n33860), .B(\key_reg[2] [2]), .C(n15489), 
         .D(n35839), .Z(key_mem_new[34])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i15069_3_lut_4_lut.init = 16'hf400;
    LUT4 i15068_3_lut_4_lut (.A(n33860), .B(\key_reg[2] [1]), .C(n15429), 
         .D(n35839), .Z(key_mem_new[33])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i15068_3_lut_4_lut.init = 16'hf400;
    LUT4 i2_2_lut_rep_264 (.A(prev_key0_reg[90]), .B(n4_adj_8438), .Z(n33568)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i2_2_lut_rep_264.init = 16'h6666;
    LUT4 i15067_3_lut_4_lut (.A(n33860), .B(\key_reg[2] [0]), .C(n15316), 
         .D(n35839), .Z(key_mem_new[32])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i15067_3_lut_4_lut.init = 16'hf400;
    LUT4 i1_3_lut_4_lut_adj_621 (.A(n33860), .B(\key_reg[3] [31]), .C(n17224), 
         .D(n35839), .Z(key_mem_new[31])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_3_lut_4_lut_adj_621.init = 16'hf400;
    LUT4 i1_3_lut_4_lut_adj_622 (.A(n33860), .B(\key_reg[3] [30]), .C(n17164), 
         .D(n35839), .Z(key_mem_new[30])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_3_lut_4_lut_adj_622.init = 16'hf400;
    LUT4 i1_3_lut_4_lut_adj_623 (.A(n33860), .B(\key_reg[3] [29]), .C(n17104), 
         .D(n35839), .Z(key_mem_new[29])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_3_lut_4_lut_adj_623.init = 16'hf400;
    LUT4 round_3__I_0_Mux_0_i11_3_lut (.A(\key_mem[12] [0]), .B(\key_mem[13] [0]), 
         .C(n33952), .Z(n11_adj_102)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_0_i11_3_lut.init = 16'hcaca;
    LUT4 i15051_2_lut_4_lut (.A(\key_reg[4] [16]), .B(n4_adj_8386), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[112])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15051_2_lut_4_lut.init = 16'hca00;
    LUT4 round_3__I_0_Mux_0_i9_3_lut (.A(\key_mem[10] [0]), .B(\key_mem[11] [0]), 
         .C(n33952), .Z(n9_adj_9102)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_0_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_0_i8_3_lut (.A(\key_mem[8] [0]), .B(\key_mem[9] [0]), 
         .C(n33952), .Z(n8_adj_9103)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_0_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_0_i5_3_lut (.A(\key_mem[6] [0]), .B(\key_mem[7] [0]), 
         .C(n33952), .Z(n5_adj_9104)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_0_i5_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_4_lut_adj_624 (.A(n33860), .B(\key_reg[3] [28]), .C(n17044), 
         .D(n35839), .Z(key_mem_new[28])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_3_lut_4_lut_adj_624.init = 16'hf400;
    LUT4 round_3__I_0_Mux_0_i4_3_lut (.A(\key_mem[4] [0]), .B(\key_mem[5] [0]), 
         .C(n33952), .Z(n4_adj_9105)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_0_i4_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_4_lut_adj_625 (.A(n33860), .B(\key_reg[3] [27]), .C(n16984), 
         .D(n35839), .Z(key_mem_new[27])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_3_lut_4_lut_adj_625.init = 16'hf400;
    LUT4 i1_3_lut_4_lut_adj_626 (.A(n33860), .B(\key_reg[3] [26]), .C(n16924), 
         .D(n35839), .Z(key_mem_new[26])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_3_lut_4_lut_adj_626.init = 16'hf400;
    LUT4 i1_3_lut_4_lut_adj_627 (.A(n33860), .B(\key_reg[3] [25]), .C(n16864), 
         .D(n35839), .Z(key_mem_new[25])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_3_lut_4_lut_adj_627.init = 16'hf400;
    LUT4 i1_3_lut_4_lut_adj_628 (.A(n33860), .B(\key_reg[3] [24]), .C(n16804), 
         .D(n35839), .Z(key_mem_new[24])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_3_lut_4_lut_adj_628.init = 16'hf400;
    LUT4 i1_3_lut_4_lut_adj_629 (.A(n33860), .B(\key_reg[3] [23]), .C(n16744), 
         .D(n35839), .Z(key_mem_new[23])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_3_lut_4_lut_adj_629.init = 16'hf400;
    LUT4 i1_3_lut_4_lut_adj_630 (.A(n33860), .B(\key_reg[3] [22]), .C(n16684), 
         .D(n35839), .Z(key_mem_new[22])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_3_lut_4_lut_adj_630.init = 16'hf400;
    LUT4 i1_3_lut_4_lut_adj_631 (.A(n33860), .B(\key_reg[3] [21]), .C(n16624), 
         .D(n35839), .Z(key_mem_new[21])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_3_lut_4_lut_adj_631.init = 16'hf400;
    LUT4 round_3__I_0_Mux_0_i2_3_lut (.A(\key_mem[2] [0]), .B(\key_mem[3] [0]), 
         .C(n33952), .Z(n2_adj_9106)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_0_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_0_i1_3_lut (.A(\key_mem[0] [0]), .B(\key_mem[1] [0]), 
         .C(n33952), .Z(n1_adj_9107)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_0_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_8_i11_3_lut (.A(\key_mem[12] [8]), .B(\key_mem[13] [8]), 
         .C(n33952), .Z(n11_adj_103)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_8_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_8_i9_3_lut (.A(\key_mem[10] [8]), .B(\key_mem[11] [8]), 
         .C(n33952), .Z(n9_adj_9109)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_8_i9_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_4_lut_adj_632 (.A(n33860), .B(\key_reg[3] [20]), .C(n16564), 
         .D(n35839), .Z(key_mem_new[20])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_3_lut_4_lut_adj_632.init = 16'hf400;
    LUT4 i1_3_lut_4_lut_adj_633 (.A(n33860), .B(\key_reg[3] [19]), .C(n16504), 
         .D(n35839), .Z(key_mem_new[19])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_3_lut_4_lut_adj_633.init = 16'hf400;
    LUT4 i1_3_lut_4_lut_adj_634 (.A(n33860), .B(\key_reg[3] [18]), .C(n16444), 
         .D(n35839), .Z(key_mem_new[18])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_3_lut_4_lut_adj_634.init = 16'hf400;
    LUT4 i1_3_lut_4_lut_adj_635 (.A(n33860), .B(\key_reg[3] [17]), .C(n16384), 
         .D(n35839), .Z(key_mem_new[17])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_3_lut_4_lut_adj_635.init = 16'hf400;
    LUT4 i1_3_lut_4_lut_adj_636 (.A(n33860), .B(\key_reg[3] [16]), .C(n16324), 
         .D(n35839), .Z(key_mem_new[16])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_3_lut_4_lut_adj_636.init = 16'hf400;
    LUT4 round_3__I_0_Mux_8_i8_3_lut (.A(\key_mem[8] [8]), .B(\key_mem[9] [8]), 
         .C(n33952), .Z(n8_adj_9110)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_8_i8_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_4_lut_adj_637 (.A(n33860), .B(\key_reg[3] [15]), .C(n16264), 
         .D(n35839), .Z(key_mem_new[15])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_3_lut_4_lut_adj_637.init = 16'hf400;
    LUT4 i1_3_lut_4_lut_adj_638 (.A(n33860), .B(\key_reg[3] [14]), .C(n16204), 
         .D(n35839), .Z(key_mem_new[14])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_3_lut_4_lut_adj_638.init = 16'hf400;
    LUT4 round_3__I_0_Mux_8_i5_3_lut (.A(\key_mem[6] [8]), .B(\key_mem[7] [8]), 
         .C(n33952), .Z(n5_adj_9111)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_8_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_8_i4_3_lut (.A(\key_mem[4] [8]), .B(\key_mem[5] [8]), 
         .C(n33952), .Z(n4_adj_9112)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_8_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_8_i2_3_lut (.A(\key_mem[2] [8]), .B(\key_mem[3] [8]), 
         .C(n33952), .Z(n2_adj_9113)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_8_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_8_i1_3_lut (.A(\key_mem[0] [8]), .B(\key_mem[1] [8]), 
         .C(n33952), .Z(n1_adj_9114)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_8_i1_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_4_lut_adj_639 (.A(n33860), .B(\key_reg[3] [13]), .C(n16144), 
         .D(n35839), .Z(key_mem_new[13])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_3_lut_4_lut_adj_639.init = 16'hf400;
    LUT4 i1_3_lut_4_lut_adj_640 (.A(n33860), .B(\key_reg[3] [12]), .C(n16084), 
         .D(n35839), .Z(key_mem_new[12])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_3_lut_4_lut_adj_640.init = 16'hf400;
    LUT4 round_3__I_0_Mux_123_i5_3_lut (.A(\key_mem[6] [123]), .B(\key_mem[7] [123]), 
         .C(n33952), .Z(n5_adj_9115)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_123_i5_3_lut.init = 16'hcaca;
    LUT4 mux_85_i91_3_lut_rep_211_4_lut (.A(prev_key0_reg[90]), .B(n4_adj_8438), 
         .C(n33859), .D(\key_reg[5] [26]), .Z(n33515)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam mux_85_i91_3_lut_rep_211_4_lut.init = 16'h6f60;
    LUT4 round_3__I_0_Mux_123_i4_3_lut (.A(\key_mem[4] [123]), .B(\key_mem[5] [123]), 
         .C(n33952), .Z(n4_adj_9116)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_123_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_7_i11_3_lut (.A(\key_mem[12] [7]), .B(\key_mem[13] [7]), 
         .C(n33952), .Z(n11_adj_104)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_7_i11_3_lut.init = 16'hcaca;
    LUT4 i15050_2_lut_4_lut (.A(\key_reg[4] [15]), .B(n4_adj_8381), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[111])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15050_2_lut_4_lut.init = 16'hca00;
    LUT4 round_3__I_0_Mux_7_i9_3_lut (.A(\key_mem[10] [7]), .B(\key_mem[11] [7]), 
         .C(n33952), .Z(n9_adj_9118)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_7_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_123_i2_3_lut (.A(\key_mem[2] [123]), .B(\key_mem[3] [123]), 
         .C(n33952), .Z(n2_adj_9119)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_123_i2_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_4_lut_adj_641 (.A(n33860), .B(\key_reg[3] [11]), .C(n16024), 
         .D(n35839), .Z(key_mem_new[11])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_3_lut_4_lut_adj_641.init = 16'hf400;
    LUT4 round_3__I_0_Mux_123_i1_3_lut (.A(\key_mem[0] [123]), .B(\key_mem[1] [123]), 
         .C(n33952), .Z(n1_adj_9120)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_123_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_7_i8_3_lut (.A(\key_mem[8] [7]), .B(\key_mem[9] [7]), 
         .C(n33952), .Z(n8_adj_9121)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_7_i8_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_4_lut_adj_642 (.A(n33860), .B(\key_reg[3] [10]), .C(n15964), 
         .D(n35839), .Z(key_mem_new[10])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_3_lut_4_lut_adj_642.init = 16'hf400;
    LUT4 i1_3_lut_4_lut_adj_643 (.A(n33860), .B(\key_reg[3] [9]), .C(n15904), 
         .D(n35839), .Z(key_mem_new[9])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_3_lut_4_lut_adj_643.init = 16'hf400;
    LUT4 i1_3_lut_4_lut_adj_644 (.A(n33860), .B(\key_reg[3] [8]), .C(n15844), 
         .D(n35839), .Z(key_mem_new[8])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_3_lut_4_lut_adj_644.init = 16'hf400;
    LUT4 i1_3_lut_4_lut_adj_645 (.A(n33860), .B(\key_reg[3] [7]), .C(n15784), 
         .D(n35839), .Z(key_mem_new[7])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_3_lut_4_lut_adj_645.init = 16'hf400;
    LUT4 i1_3_lut_4_lut_adj_646 (.A(n33860), .B(\key_reg[3] [6]), .C(n15724), 
         .D(n35839), .Z(key_mem_new[6])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_3_lut_4_lut_adj_646.init = 16'hf400;
    LUT4 i1_3_lut_4_lut_adj_647 (.A(n33860), .B(\key_reg[3] [5]), .C(n15664), 
         .D(n35839), .Z(key_mem_new[5])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_3_lut_4_lut_adj_647.init = 16'hf400;
    LUT4 i1_3_lut_4_lut_adj_648 (.A(n33860), .B(\key_reg[3] [4]), .C(n15604), 
         .D(n35839), .Z(key_mem_new[4])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_3_lut_4_lut_adj_648.init = 16'hf400;
    LUT4 i1_3_lut_4_lut_adj_649 (.A(n33860), .B(\key_reg[3] [3]), .C(n15544), 
         .D(n35839), .Z(key_mem_new[3])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_3_lut_4_lut_adj_649.init = 16'hf400;
    LUT4 i1_3_lut_4_lut_adj_650 (.A(n33860), .B(\key_reg[3] [2]), .C(n15484), 
         .D(n35839), .Z(key_mem_new[2])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_3_lut_4_lut_adj_650.init = 16'hf400;
    LUT4 i1_3_lut_4_lut_adj_651 (.A(n33860), .B(\key_reg[3] [1]), .C(n15424), 
         .D(n35839), .Z(key_mem_new[1])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_3_lut_4_lut_adj_651.init = 16'hf400;
    LUT4 round_3__I_0_Mux_122_i11_3_lut (.A(\key_mem[12] [122]), .B(\key_mem[13] [122]), 
         .C(n33952), .Z(n11_adj_105)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_122_i11_3_lut.init = 16'hcaca;
    LUT4 mux_9_i65_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [64]), 
         .D(key_mem_new[64]), .Z(key_mem_0__127__N_6752[64])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i65_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i40_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [39]), 
         .D(key_mem_new[39]), .Z(key_mem_0__127__N_6752[39])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i40_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i41_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [40]), 
         .D(key_mem_new[40]), .Z(key_mem_0__127__N_6752[40])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i41_3_lut_4_lut.init = 16'hf4b0;
    LUT4 round_3__I_0_Mux_7_i5_3_lut (.A(\key_mem[6] [7]), .B(\key_mem[7] [7]), 
         .C(n33952), .Z(n5_adj_9123)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_7_i5_3_lut.init = 16'hcaca;
    LUT4 mux_9_i42_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [41]), 
         .D(key_mem_new[41]), .Z(key_mem_0__127__N_6752[41])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i42_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i43_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [42]), 
         .D(key_mem_new[42]), .Z(key_mem_0__127__N_6752[42])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i43_3_lut_4_lut.init = 16'hf4b0;
    LUT4 round_3__I_0_Mux_122_i9_3_lut (.A(\key_mem[10] [122]), .B(\key_mem[11] [122]), 
         .C(n33952), .Z(n9_adj_9124)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_122_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_7_i4_3_lut (.A(\key_mem[4] [7]), .B(\key_mem[5] [7]), 
         .C(n33952), .Z(n4_adj_9125)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_7_i4_3_lut.init = 16'hcaca;
    LUT4 mux_9_i44_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [43]), 
         .D(key_mem_new[43]), .Z(key_mem_0__127__N_6752[43])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i44_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i45_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [44]), 
         .D(key_mem_new[44]), .Z(key_mem_0__127__N_6752[44])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i45_3_lut_4_lut.init = 16'hf4b0;
    LUT4 round_3__I_0_Mux_7_i2_3_lut (.A(\key_mem[2] [7]), .B(\key_mem[3] [7]), 
         .C(n33952), .Z(n2_adj_9126)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_7_i2_3_lut.init = 16'hcaca;
    LUT4 mux_9_i46_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [45]), 
         .D(key_mem_new[45]), .Z(key_mem_0__127__N_6752[45])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i46_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i47_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [46]), 
         .D(key_mem_new[46]), .Z(key_mem_0__127__N_6752[46])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i47_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i48_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [47]), 
         .D(key_mem_new[47]), .Z(key_mem_0__127__N_6752[47])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i48_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i49_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [48]), 
         .D(key_mem_new[48]), .Z(key_mem_0__127__N_6752[48])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i49_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i50_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [49]), 
         .D(key_mem_new[49]), .Z(key_mem_0__127__N_6752[49])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i50_3_lut_4_lut.init = 16'hf4b0;
    LUT4 round_3__I_0_Mux_122_i8_3_lut (.A(\key_mem[8] [122]), .B(\key_mem[9] [122]), 
         .C(n33952), .Z(n8_adj_9127)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_122_i8_3_lut.init = 16'hcaca;
    LUT4 mux_9_i51_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [50]), 
         .D(key_mem_new[50]), .Z(key_mem_0__127__N_6752[50])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i51_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i52_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [51]), 
         .D(key_mem_new[51]), .Z(key_mem_0__127__N_6752[51])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i52_3_lut_4_lut.init = 16'hf4b0;
    LUT4 round_3__I_0_Mux_7_i1_3_lut (.A(\key_mem[0] [7]), .B(\key_mem[1] [7]), 
         .C(n33952), .Z(n1_adj_9128)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_7_i1_3_lut.init = 16'hcaca;
    LUT4 mux_9_i53_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [52]), 
         .D(key_mem_new[52]), .Z(key_mem_0__127__N_6752[52])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i53_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i54_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [53]), 
         .D(key_mem_new[53]), .Z(key_mem_0__127__N_6752[53])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i54_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i55_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [54]), 
         .D(key_mem_new[54]), .Z(key_mem_0__127__N_6752[54])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i55_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i56_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [55]), 
         .D(key_mem_new[55]), .Z(key_mem_0__127__N_6752[55])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i56_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i57_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [56]), 
         .D(key_mem_new[56]), .Z(key_mem_0__127__N_6752[56])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i57_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i58_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [57]), 
         .D(key_mem_new[57]), .Z(key_mem_0__127__N_6752[57])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i58_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i59_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [58]), 
         .D(key_mem_new[58]), .Z(key_mem_0__127__N_6752[58])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i59_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i60_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [59]), 
         .D(key_mem_new[59]), .Z(key_mem_0__127__N_6752[59])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i60_3_lut_4_lut.init = 16'hf4b0;
    LUT4 round_3__I_0_Mux_122_i5_3_lut (.A(\key_mem[6] [122]), .B(\key_mem[7] [122]), 
         .C(n33952), .Z(n5_adj_9129)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_122_i5_3_lut.init = 16'hcaca;
    LUT4 i6_2_lut_3_lut_adj_652 (.A(prev_key1_reg[58]), .B(n33618), .C(keymem_sboxw[26]), 
         .Z(n16917)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;
    defparam i6_2_lut_3_lut_adj_652.init = 16'h9696;
    LUT4 round_3__I_0_Mux_26_i11_3_lut (.A(\key_mem[12] [26]), .B(\key_mem[13] [26]), 
         .C(n33952), .Z(n11_adj_106)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_26_i11_3_lut.init = 16'hcaca;
    LUT4 i15049_2_lut_4_lut (.A(\key_reg[4] [14]), .B(n4_adj_8377), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[110])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15049_2_lut_4_lut.init = 16'hca00;
    LUT4 round_3__I_0_Mux_26_i9_3_lut (.A(\key_mem[10] [26]), .B(\key_mem[11] [26]), 
         .C(n33952), .Z(n9_adj_9131)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_26_i9_3_lut.init = 16'hcaca;
    LUT4 mux_9_i61_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [60]), 
         .D(key_mem_new[60]), .Z(key_mem_0__127__N_6752[60])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i61_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i62_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [61]), 
         .D(key_mem_new[61]), .Z(key_mem_0__127__N_6752[61])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i62_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i63_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [62]), 
         .D(key_mem_new[62]), .Z(key_mem_0__127__N_6752[62])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i63_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i64_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [63]), 
         .D(key_mem_new[63]), .Z(key_mem_0__127__N_6752[63])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i64_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i1_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [0]), 
         .D(key_mem_new[0]), .Z(key_mem_0__127__N_6752[0])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i1_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i2_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [1]), 
         .D(key_mem_new[1]), .Z(key_mem_0__127__N_6752[1])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i2_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i3_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [2]), 
         .D(key_mem_new[2]), .Z(key_mem_0__127__N_6752[2])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i3_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i4_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [3]), 
         .D(key_mem_new[3]), .Z(key_mem_0__127__N_6752[3])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i4_3_lut_4_lut.init = 16'hf4b0;
    LUT4 round_3__I_0_Mux_26_i8_3_lut (.A(\key_mem[8] [26]), .B(\key_mem[9] [26]), 
         .C(n33952), .Z(n8_adj_9132)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_26_i8_3_lut.init = 16'hcaca;
    LUT4 mux_9_i5_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [4]), 
         .D(key_mem_new[4]), .Z(key_mem_0__127__N_6752[4])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i5_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i6_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [5]), 
         .D(key_mem_new[5]), .Z(key_mem_0__127__N_6752[5])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i6_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i7_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [6]), 
         .D(key_mem_new[6]), .Z(key_mem_0__127__N_6752[6])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i7_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i8_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [7]), 
         .D(key_mem_new[7]), .Z(key_mem_0__127__N_6752[7])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i8_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i9_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [8]), 
         .D(key_mem_new[8]), .Z(key_mem_0__127__N_6752[8])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i9_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i10_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [9]), 
         .D(key_mem_new[9]), .Z(key_mem_0__127__N_6752[9])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i10_3_lut_4_lut.init = 16'hf4b0;
    LUT4 round_3__I_0_Mux_26_i5_3_lut (.A(\key_mem[6] [26]), .B(\key_mem[7] [26]), 
         .C(n33952), .Z(n5_adj_9133)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_26_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_26_i4_3_lut (.A(\key_mem[4] [26]), .B(\key_mem[5] [26]), 
         .C(n33952), .Z(n4_adj_9134)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_26_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_26_i2_3_lut (.A(\key_mem[2] [26]), .B(\key_mem[3] [26]), 
         .C(n33952), .Z(n2_adj_9135)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_26_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_26_i1_3_lut (.A(\key_mem[0] [26]), .B(\key_mem[1] [26]), 
         .C(n33952), .Z(n1_adj_9136)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_26_i1_3_lut.init = 16'hcaca;
    LUT4 mux_9_i11_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [10]), 
         .D(key_mem_new[10]), .Z(key_mem_0__127__N_6752[10])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i11_3_lut_4_lut.init = 16'hf4b0;
    LUT4 round_3__I_0_Mux_122_i4_3_lut (.A(\key_mem[4] [122]), .B(\key_mem[5] [122]), 
         .C(n33952), .Z(n4_adj_9137)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_122_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_6_i11_3_lut (.A(\key_mem[12] [6]), .B(\key_mem[13] [6]), 
         .C(n33952), .Z(n11_adj_107)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_6_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_6_i9_3_lut (.A(\key_mem[10] [6]), .B(\key_mem[11] [6]), 
         .C(n33952), .Z(n9_adj_9139)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_6_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_6_i8_3_lut (.A(\key_mem[8] [6]), .B(\key_mem[9] [6]), 
         .C(n33952), .Z(n8_adj_9140)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_6_i8_3_lut.init = 16'hcaca;
    LUT4 mux_9_i12_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [11]), 
         .D(key_mem_new[11]), .Z(key_mem_0__127__N_6752[11])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i12_3_lut_4_lut.init = 16'hf4b0;
    LUT4 round_3__I_0_Mux_6_i5_3_lut (.A(\key_mem[6] [6]), .B(\key_mem[7] [6]), 
         .C(n33952), .Z(n5_adj_9141)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_6_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_6_i4_3_lut (.A(\key_mem[4] [6]), .B(\key_mem[5] [6]), 
         .C(n33952), .Z(n4_adj_9142)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_6_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_6_i2_3_lut (.A(\key_mem[2] [6]), .B(\key_mem[3] [6]), 
         .C(n33952), .Z(n2_adj_9143)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_6_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_6_i1_3_lut (.A(\key_mem[0] [6]), .B(\key_mem[1] [6]), 
         .C(n33952), .Z(n1_adj_9144)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_6_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_122_i2_3_lut (.A(\key_mem[2] [122]), .B(\key_mem[3] [122]), 
         .C(n33952), .Z(n2_adj_9145)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_122_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_5_i11_3_lut (.A(\key_mem[12] [5]), .B(\key_mem[13] [5]), 
         .C(n33952), .Z(n11_adj_108)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_5_i11_3_lut.init = 16'hcaca;
    LUT4 i15048_2_lut_4_lut (.A(\key_reg[4] [13]), .B(n4_adj_8373), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[109])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15048_2_lut_4_lut.init = 16'hca00;
    LUT4 mux_9_i13_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [12]), 
         .D(key_mem_new[12]), .Z(key_mem_0__127__N_6752[12])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i13_3_lut_4_lut.init = 16'hf4b0;
    LUT4 round_3__I_0_Mux_5_i9_3_lut (.A(\key_mem[10] [5]), .B(\key_mem[11] [5]), 
         .C(n33952), .Z(n9_adj_9147)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_5_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_5_i8_3_lut (.A(\key_mem[8] [5]), .B(\key_mem[9] [5]), 
         .C(n33952), .Z(n8_adj_9148)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_5_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_5_i5_3_lut (.A(\key_mem[6] [5]), .B(\key_mem[7] [5]), 
         .C(n33952), .Z(n5_adj_9149)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_5_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_5_i4_3_lut (.A(\key_mem[4] [5]), .B(\key_mem[5] [5]), 
         .C(n33952), .Z(n4_adj_9150)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_5_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_122_i1_3_lut (.A(\key_mem[0] [122]), .B(\key_mem[1] [122]), 
         .C(n33952), .Z(n1_adj_9151)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_122_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_5_i2_3_lut (.A(\key_mem[2] [5]), .B(\key_mem[3] [5]), 
         .C(n33952), .Z(n2_adj_9152)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_5_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_5_i1_3_lut (.A(\key_mem[0] [5]), .B(\key_mem[1] [5]), 
         .C(n33952), .Z(n1_adj_9153)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_5_i1_3_lut.init = 16'hcaca;
    LUT4 mux_9_i14_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [13]), 
         .D(key_mem_new[13]), .Z(key_mem_0__127__N_6752[13])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i14_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i2_2_lut_rep_267 (.A(prev_key0_reg[89]), .B(n4_adj_8430), .Z(n33571)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i2_2_lut_rep_267.init = 16'h6666;
    LUT4 round_3__I_0_Mux_4_i11_3_lut (.A(\key_mem[12] [4]), .B(\key_mem[13] [4]), 
         .C(n33952), .Z(n11_adj_109)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_4_i11_3_lut.init = 16'hcaca;
    LUT4 mux_9_i15_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [14]), 
         .D(key_mem_new[14]), .Z(key_mem_0__127__N_6752[14])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i15_3_lut_4_lut.init = 16'hf4b0;
    LUT4 round_3__I_0_Mux_121_i11_3_lut (.A(\key_mem[12] [121]), .B(\key_mem[13] [121]), 
         .C(n33952), .Z(n11_adj_110)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_121_i11_3_lut.init = 16'hcaca;
    LUT4 mux_9_i16_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [15]), 
         .D(key_mem_new[15]), .Z(key_mem_0__127__N_6752[15])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i16_3_lut_4_lut.init = 16'hf4b0;
    LUT4 round_3__I_0_Mux_4_i9_3_lut (.A(\key_mem[10] [4]), .B(\key_mem[11] [4]), 
         .C(n33952), .Z(n9_adj_9156)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_4_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_4_i8_3_lut (.A(\key_mem[8] [4]), .B(\key_mem[9] [4]), 
         .C(n33952), .Z(n8_adj_9157)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_4_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_4_i5_3_lut (.A(\key_mem[6] [4]), .B(\key_mem[7] [4]), 
         .C(n33952), .Z(n5_adj_9158)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_4_i5_3_lut.init = 16'hcaca;
    LUT4 i15047_2_lut_4_lut (.A(\key_reg[4] [12]), .B(n4_adj_8367), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[108])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15047_2_lut_4_lut.init = 16'hca00;
    LUT4 round_3__I_0_Mux_4_i4_3_lut (.A(\key_mem[4] [4]), .B(\key_mem[5] [4]), 
         .C(n33952), .Z(n4_adj_9159)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_4_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_4_i2_3_lut (.A(\key_mem[2] [4]), .B(\key_mem[3] [4]), 
         .C(n33952), .Z(n2_adj_9160)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_4_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_4_i1_3_lut (.A(\key_mem[0] [4]), .B(\key_mem[1] [4]), 
         .C(n33952), .Z(n1_adj_9161)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_4_i1_3_lut.init = 16'hcaca;
    LUT4 mux_85_i90_3_lut_rep_212_4_lut (.A(prev_key0_reg[89]), .B(n4_adj_8430), 
         .C(n33859), .D(\key_reg[5] [25]), .Z(n33516)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam mux_85_i90_3_lut_rep_212_4_lut.init = 16'h6f60;
    LUT4 round_3__I_0_Mux_3_i11_3_lut (.A(\key_mem[12] [3]), .B(\key_mem[13] [3]), 
         .C(n33952), .Z(n11_adj_111)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_3_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_121_i9_3_lut (.A(\key_mem[10] [121]), .B(\key_mem[11] [121]), 
         .C(n33952), .Z(n9_adj_9163)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_121_i9_3_lut.init = 16'hcaca;
    LUT4 mux_9_i17_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [16]), 
         .D(key_mem_new[16]), .Z(key_mem_0__127__N_6752[16])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i17_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i18_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [17]), 
         .D(key_mem_new[17]), .Z(key_mem_0__127__N_6752[17])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i18_3_lut_4_lut.init = 16'hf4b0;
    LUT4 round_3__I_0_Mux_3_i9_3_lut (.A(\key_mem[10] [3]), .B(\key_mem[11] [3]), 
         .C(n33952), .Z(n9_adj_9164)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_3_i9_3_lut.init = 16'hcaca;
    LUT4 mux_9_i19_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [18]), 
         .D(key_mem_new[18]), .Z(key_mem_0__127__N_6752[18])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i19_3_lut_4_lut.init = 16'hf4b0;
    LUT4 round_3__I_0_Mux_3_i8_3_lut (.A(\key_mem[8] [3]), .B(\key_mem[9] [3]), 
         .C(n33952), .Z(n8_adj_9165)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_3_i8_3_lut.init = 16'hcaca;
    LUT4 mux_9_i20_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [19]), 
         .D(key_mem_new[19]), .Z(key_mem_0__127__N_6752[19])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i20_3_lut_4_lut.init = 16'hf4b0;
    L6MUX21 i25244 (.D0(n30399), .D1(n30400), .SD(\muxed_round_nr[2] ), 
            .Z(n30403));
    L6MUX21 i25245 (.D0(n30401), .D1(n33394), .SD(\muxed_round_nr[2] ), 
            .Z(n30404));
    LUT4 round_3__I_0_Mux_3_i5_3_lut (.A(\key_mem[6] [3]), .B(\key_mem[7] [3]), 
         .C(n33952), .Z(n5_adj_9166)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_3_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_3_i4_3_lut (.A(\key_mem[4] [3]), .B(\key_mem[5] [3]), 
         .C(n33952), .Z(n4_adj_9167)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_3_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_105_i2_3_lut (.A(\key_mem[2] [105]), .B(\key_mem[3] [105]), 
         .C(n33952), .Z(n2)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_105_i2_3_lut.init = 16'hcaca;
    LUT4 mux_9_i21_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [20]), 
         .D(key_mem_new[20]), .Z(key_mem_0__127__N_6752[20])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i21_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i22_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [21]), 
         .D(key_mem_new[21]), .Z(key_mem_0__127__N_6752[21])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i22_3_lut_4_lut.init = 16'hf4b0;
    LUT4 round_3__I_0_Mux_3_i2_3_lut (.A(\key_mem[2] [3]), .B(\key_mem[3] [3]), 
         .C(n33952), .Z(n2_adj_9168)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_3_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_3_i1_3_lut (.A(\key_mem[0] [3]), .B(\key_mem[1] [3]), 
         .C(n33952), .Z(n1_adj_9169)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_3_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_2_i11_3_lut (.A(\key_mem[12] [2]), .B(\key_mem[13] [2]), 
         .C(n33952), .Z(n11_adj_112)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_2_i11_3_lut.init = 16'hcaca;
    LUT4 i15046_2_lut_4_lut (.A(\key_reg[4] [11]), .B(n4_adj_8361), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[107])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15046_2_lut_4_lut.init = 16'hca00;
    LUT4 round_3__I_0_Mux_2_i9_3_lut (.A(\key_mem[10] [2]), .B(\key_mem[11] [2]), 
         .C(n33952), .Z(n9_adj_9171)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_2_i9_3_lut.init = 16'hcaca;
    L6MUX21 i25251 (.D0(n30406), .D1(n30407), .SD(\muxed_round_nr[2] ), 
            .Z(n30410));
    FD1P3IX prev_key0_reg__i1 (.D(prev_key0_new_127__N_4659[1]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[1])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i1.GSR = "DISABLED";
    L6MUX21 i25252 (.D0(n30408), .D1(n33396), .SD(\muxed_round_nr[2] ), 
            .Z(n30411));
    LUT4 round_3__I_0_Mux_2_i8_3_lut (.A(\key_mem[8] [2]), .B(\key_mem[9] [2]), 
         .C(n33952), .Z(n8_adj_9172)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_2_i8_3_lut.init = 16'hcaca;
    L6MUX21 i25258 (.D0(n30413), .D1(n30414), .SD(\muxed_round_nr[2] ), 
            .Z(n30417));
    LUT4 round_3__I_0_Mux_2_i5_3_lut (.A(\key_mem[6] [2]), .B(\key_mem[7] [2]), 
         .C(n33952), .Z(n5_adj_9173)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_2_i5_3_lut.init = 16'hcaca;
    L6MUX21 i25259 (.D0(n30415), .D1(n33397), .SD(\muxed_round_nr[2] ), 
            .Z(n30418));
    LUT4 round_3__I_0_Mux_2_i4_3_lut (.A(\key_mem[4] [2]), .B(\key_mem[5] [2]), 
         .C(n33952), .Z(n4_adj_9174)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_2_i4_3_lut.init = 16'hcaca;
    L6MUX21 i25265 (.D0(n30420), .D1(n30421), .SD(\muxed_round_nr[2] ), 
            .Z(n30424));
    LUT4 round_3__I_0_Mux_2_i2_3_lut (.A(\key_mem[2] [2]), .B(\key_mem[3] [2]), 
         .C(n33952), .Z(n2_adj_9175)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_2_i2_3_lut.init = 16'hcaca;
    L6MUX21 i25266 (.D0(n30422), .D1(n33399), .SD(\muxed_round_nr[2] ), 
            .Z(n30425));
    LUT4 round_3__I_0_Mux_2_i1_3_lut (.A(\key_mem[0] [2]), .B(\key_mem[1] [2]), 
         .C(n33952), .Z(n1_adj_9176)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_2_i1_3_lut.init = 16'hcaca;
    L6MUX21 i25272 (.D0(n30427), .D1(n30428), .SD(\muxed_round_nr[2] ), 
            .Z(n30431));
    LUT4 mux_9_i23_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [22]), 
         .D(key_mem_new[22]), .Z(key_mem_0__127__N_6752[22])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i23_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i6_2_lut_3_lut_adj_653 (.A(prev_key1_reg[56]), .B(n33619), .C(keymem_sboxw[24]), 
         .Z(n16797)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;
    defparam i6_2_lut_3_lut_adj_653.init = 16'h9696;
    L6MUX21 i25273 (.D0(n30429), .D1(n33401), .SD(\muxed_round_nr[2] ), 
            .Z(n30432));
    LUT4 round_3__I_0_Mux_1_i11_3_lut (.A(\key_mem[12] [1]), .B(\key_mem[13] [1]), 
         .C(n33952), .Z(n11_adj_113)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_1_i11_3_lut.init = 16'hcaca;
    L6MUX21 i25279 (.D0(n30434), .D1(n30435), .SD(\muxed_round_nr[2] ), 
            .Z(n30438));
    LUT4 mux_9_i24_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [23]), 
         .D(key_mem_new[23]), .Z(key_mem_0__127__N_6752[23])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i24_3_lut_4_lut.init = 16'hf4b0;
    L6MUX21 i25280 (.D0(n30436), .D1(n33403), .SD(\muxed_round_nr[2] ), 
            .Z(n30439));
    LUT4 mux_9_i25_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [24]), 
         .D(key_mem_new[24]), .Z(key_mem_0__127__N_6752[24])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i25_3_lut_4_lut.init = 16'hf4b0;
    L6MUX21 i25286 (.D0(n30441), .D1(n30442), .SD(\muxed_round_nr[2] ), 
            .Z(n30445));
    LUT4 round_3__I_0_Mux_1_i9_3_lut (.A(\key_mem[10] [1]), .B(\key_mem[11] [1]), 
         .C(n33952), .Z(n9_adj_9178)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_1_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_1_i8_3_lut (.A(\key_mem[8] [1]), .B(\key_mem[9] [1]), 
         .C(n33952), .Z(n8_adj_9179)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_1_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_1_i5_3_lut (.A(\key_mem[6] [1]), .B(\key_mem[7] [1]), 
         .C(n33952), .Z(n5_adj_9180)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_1_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_1_i4_3_lut (.A(\key_mem[4] [1]), .B(\key_mem[5] [1]), 
         .C(n33952), .Z(n4_adj_9181)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_1_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_1_i2_3_lut (.A(\key_mem[2] [1]), .B(\key_mem[3] [1]), 
         .C(n33952), .Z(n2_adj_9182)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_1_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_1_i1_3_lut (.A(\key_mem[0] [1]), .B(\key_mem[1] [1]), 
         .C(n33952), .Z(n1_adj_9183)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_1_i1_3_lut.init = 16'hcaca;
    LUT4 i2_2_lut_rep_269 (.A(prev_key0_reg[88]), .B(n4_adj_8428), .Z(n33573)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i2_2_lut_rep_269.init = 16'h6666;
    LUT4 round_3__I_0_Mux_46_i11_3_lut (.A(\key_mem[12] [46]), .B(\key_mem[13] [46]), 
         .C(n33952), .Z(n11_adj_114)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_46_i11_3_lut.init = 16'hcaca;
    LUT4 i15045_2_lut_4_lut (.A(\key_reg[4] [10]), .B(n4), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[106])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15045_2_lut_4_lut.init = 16'hca00;
    LUT4 round_3__I_0_Mux_46_i9_3_lut (.A(\key_mem[10] [46]), .B(\key_mem[11] [46]), 
         .C(n33952), .Z(n9_adj_9185)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_46_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_46_i8_3_lut (.A(\key_mem[8] [46]), .B(\key_mem[9] [46]), 
         .C(n33952), .Z(n8_adj_9186)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_46_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_46_i5_3_lut (.A(\key_mem[6] [46]), .B(\key_mem[7] [46]), 
         .C(n33952), .Z(n5_adj_9187)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_46_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_46_i4_3_lut (.A(\key_mem[4] [46]), .B(\key_mem[5] [46]), 
         .C(n33952), .Z(n4_adj_9188)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_46_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_46_i2_3_lut (.A(\key_mem[2] [46]), .B(\key_mem[3] [46]), 
         .C(n33952), .Z(n2_adj_9189)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_46_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_46_i1_3_lut (.A(\key_mem[0] [46]), .B(\key_mem[1] [46]), 
         .C(maxfan_replicated_net_23), .Z(n1_adj_9190)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_46_i1_3_lut.init = 16'hcaca;
    LUT4 mux_85_i89_3_lut_rep_213_4_lut (.A(prev_key0_reg[88]), .B(n4_adj_8428), 
         .C(n33859), .D(\key_reg[5] [24]), .Z(n33517)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam mux_85_i89_3_lut_rep_213_4_lut.init = 16'h6f60;
    LUT4 round_3__I_0_Mux_45_i11_3_lut (.A(\key_mem[12] [45]), .B(\key_mem[13] [45]), 
         .C(maxfan_replicated_net_23), .Z(n11_adj_115)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_45_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_45_i9_3_lut (.A(\key_mem[10] [45]), .B(\key_mem[11] [45]), 
         .C(maxfan_replicated_net_23), .Z(n9_adj_9192)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_45_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_45_i8_3_lut (.A(\key_mem[8] [45]), .B(\key_mem[9] [45]), 
         .C(maxfan_replicated_net_23), .Z(n8_adj_9193)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_45_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_45_i5_3_lut (.A(\key_mem[6] [45]), .B(\key_mem[7] [45]), 
         .C(maxfan_replicated_net_23), .Z(n5_adj_9194)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_45_i5_3_lut.init = 16'hcaca;
    FD1P3IX prev_key0_reg__i2 (.D(prev_key0_new_127__N_4659[2]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[2])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i2.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i3 (.D(prev_key0_new_127__N_4659[3]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[3])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i3.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i4 (.D(prev_key0_new_127__N_4659[4]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[4])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i4.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i5 (.D(prev_key0_new_127__N_4659[5]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[5])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i5.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i6 (.D(prev_key0_new_127__N_4659[6]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[6])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i6.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i7 (.D(prev_key0_new_127__N_4659[7]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[7])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i7.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i8 (.D(prev_key0_new_127__N_4659[8]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[8])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i8.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i9 (.D(prev_key0_new_127__N_4659[9]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[9])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i9.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i10 (.D(prev_key0_new_127__N_4659[10]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[10])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i10.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i11 (.D(prev_key0_new_127__N_4659[11]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[11])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i11.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i12 (.D(prev_key0_new_127__N_4659[12]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[12])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i12.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i13 (.D(prev_key0_new_127__N_4659[13]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[13])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i13.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i14 (.D(prev_key0_new_127__N_4659[14]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[14])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i14.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i15 (.D(prev_key0_new_127__N_4659[15]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[15])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i15.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i16 (.D(prev_key0_new_127__N_4659[16]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[16])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i16.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i17 (.D(prev_key0_new_127__N_4659[17]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[17])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i17.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i18 (.D(prev_key0_new_127__N_4659[18]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[18])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i18.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i19 (.D(prev_key0_new_127__N_4659[19]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[19])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i19.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i20 (.D(prev_key0_new_127__N_4659[20]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[20])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i20.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i21 (.D(prev_key0_new_127__N_4659[21]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[21])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i21.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i22 (.D(prev_key0_new_127__N_4659[22]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[22])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i22.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i23 (.D(prev_key0_new_127__N_4659[23]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[23])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i23.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i24 (.D(prev_key0_new_127__N_4659[24]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[24])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i24.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i25 (.D(prev_key0_new_127__N_4659[25]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[25])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i25.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i26 (.D(prev_key0_new_127__N_4659[26]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[26])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i26.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i27 (.D(prev_key0_new_127__N_4659[27]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[27])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i27.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i28 (.D(prev_key0_new_127__N_4659[28]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[28])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i28.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i29 (.D(prev_key0_new_127__N_4659[29]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[29])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i29.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i30 (.D(prev_key0_new_127__N_4659[30]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[30])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i30.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i31 (.D(prev_key0_new_127__N_4659[31]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[31])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i31.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i32 (.D(prev_key0_new_127__N_4659[32]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[32])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i32.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i33 (.D(prev_key0_new_127__N_4659[33]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[33])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i33.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i34 (.D(prev_key0_new_127__N_4659[34]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[34])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i34.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i35 (.D(prev_key0_new_127__N_4659[35]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[35])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i35.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i36 (.D(prev_key0_new_127__N_4659[36]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[36])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i36.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i37 (.D(prev_key0_new_127__N_4659[37]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[37])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i37.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i38 (.D(prev_key0_new_127__N_4659[38]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[38])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i38.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i39 (.D(prev_key0_new_127__N_4659[39]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[39])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i39.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i40 (.D(prev_key0_new_127__N_4659[40]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[40])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i40.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i41 (.D(prev_key0_new_127__N_4659[41]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[41])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i41.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i42 (.D(prev_key0_new_127__N_4659[42]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[42])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i42.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i43 (.D(prev_key0_new_127__N_4659[43]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[43])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i43.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i44 (.D(prev_key0_new_127__N_4659[44]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[44])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i44.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i45 (.D(prev_key0_new_127__N_4659[45]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[45])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i45.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i46 (.D(prev_key0_new_127__N_4659[46]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[46])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i46.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i47 (.D(prev_key0_new_127__N_4659[47]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[47])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i47.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i48 (.D(prev_key0_new_127__N_4659[48]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[48])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i48.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i49 (.D(prev_key0_new_127__N_4659[49]), .SP(clk_c_enable_54), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[49])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i49.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i50 (.D(prev_key0_new_127__N_4659[50]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[50])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i50.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i51 (.D(prev_key0_new_127__N_4659[51]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[51])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i51.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i52 (.D(prev_key0_new_127__N_4659[52]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[52])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i52.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i53 (.D(prev_key0_new_127__N_4659[53]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[53])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i53.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i54 (.D(prev_key0_new_127__N_4659[54]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[54])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i54.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i55 (.D(prev_key0_new_127__N_4659[55]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[55])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i55.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i56 (.D(prev_key0_new_127__N_4659[56]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[56])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i56.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i57 (.D(prev_key0_new_127__N_4659[57]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[57])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i57.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i58 (.D(prev_key0_new_127__N_4659[58]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[58])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i58.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i59 (.D(prev_key0_new_127__N_4659[59]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[59])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i59.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i60 (.D(prev_key0_new_127__N_4659[60]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[60])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i60.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i61 (.D(prev_key0_new_127__N_4659[61]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[61])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i61.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i62 (.D(prev_key0_new_127__N_4659[62]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[62])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i62.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i63 (.D(prev_key0_new_127__N_4659[63]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[63])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i63.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i64 (.D(prev_key0_new_127__N_4659[64]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[64])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i64.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i65 (.D(prev_key0_new_127__N_4659[65]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[65])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i65.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i66 (.D(prev_key0_new_127__N_4659[66]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[66])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i66.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i67 (.D(prev_key0_new_127__N_4659[67]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[67])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i67.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i68 (.D(prev_key0_new_127__N_4659[68]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[68])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i68.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i69 (.D(prev_key0_new_127__N_4659[69]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[69])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i69.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i70 (.D(prev_key0_new_127__N_4659[70]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[70])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i70.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i71 (.D(prev_key0_new_127__N_4659[71]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[71])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i71.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i72 (.D(prev_key0_new_127__N_4659[72]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[72])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i72.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i73 (.D(prev_key0_new_127__N_4659[73]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[73])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i73.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i74 (.D(prev_key0_new_127__N_4659[74]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[74])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i74.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i75 (.D(prev_key0_new_127__N_4659[75]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[75])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i75.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i76 (.D(prev_key0_new_127__N_4659[76]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[76])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i76.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i77 (.D(prev_key0_new_127__N_4659[77]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[77])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i77.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i78 (.D(prev_key0_new_127__N_4659[78]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[78])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i78.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i79 (.D(prev_key0_new_127__N_4659[79]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[79])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i79.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i80 (.D(prev_key0_new_127__N_4659[80]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[80])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i80.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i81 (.D(prev_key0_new_127__N_4659[81]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[81])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i81.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i82 (.D(prev_key0_new_127__N_4659[82]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[82])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i82.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i83 (.D(prev_key0_new_127__N_4659[83]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[83])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i83.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i84 (.D(prev_key0_new_127__N_4659[84]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[84])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i84.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i85 (.D(prev_key0_new_127__N_4659[85]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[85])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i85.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i86 (.D(prev_key0_new_127__N_4659[86]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[86])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i86.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i87 (.D(prev_key0_new_127__N_4659[87]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[87])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i87.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i88 (.D(prev_key0_new_127__N_4659[88]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[88])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i88.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i89 (.D(prev_key0_new_127__N_4659[89]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[89])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i89.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i90 (.D(prev_key0_new_127__N_4659[90]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[90])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i90.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i91 (.D(prev_key0_new_127__N_4659[91]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[91])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i91.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i92 (.D(prev_key0_new_127__N_4659[92]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[92])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i92.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i93 (.D(prev_key0_new_127__N_4659[93]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[93])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i93.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i94 (.D(prev_key0_new_127__N_4659[94]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[94])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i94.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i95 (.D(prev_key0_new_127__N_4659[95]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[95])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i95.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i96 (.D(prev_key0_new_127__N_4659[96]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[96])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i96.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i97 (.D(prev_key0_new_127__N_4659[97]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[97])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i97.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i98 (.D(prev_key0_new_127__N_4659[98]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[98])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i98.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i99 (.D(prev_key0_new_127__N_4659[99]), .SP(clk_c_enable_104), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[99])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i99.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i100 (.D(prev_key0_new_127__N_4659[100]), .SP(clk_c_enable_132), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[100])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i100.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i101 (.D(prev_key0_new_127__N_4659[101]), .SP(clk_c_enable_132), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[101])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i101.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i102 (.D(prev_key0_new_127__N_4659[102]), .SP(clk_c_enable_132), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[102])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i102.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i103 (.D(prev_key0_new_127__N_4659[103]), .SP(clk_c_enable_132), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[103])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i103.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i104 (.D(prev_key0_new_127__N_4659[104]), .SP(clk_c_enable_132), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[104])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i104.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i105 (.D(prev_key0_new_127__N_4659[105]), .SP(clk_c_enable_132), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[105])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i105.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i106 (.D(prev_key0_new_127__N_4659[106]), .SP(clk_c_enable_132), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[106])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i106.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i107 (.D(prev_key0_new_127__N_4659[107]), .SP(clk_c_enable_132), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[107])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i107.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i108 (.D(prev_key0_new_127__N_4659[108]), .SP(clk_c_enable_132), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[108])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i108.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i109 (.D(prev_key0_new_127__N_4659[109]), .SP(clk_c_enable_132), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[109])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i109.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i110 (.D(prev_key0_new_127__N_4659[110]), .SP(clk_c_enable_132), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[110])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i110.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i111 (.D(prev_key0_new_127__N_4659[111]), .SP(clk_c_enable_132), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[111])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i111.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i112 (.D(prev_key0_new_127__N_4659[112]), .SP(clk_c_enable_132), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[112])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i112.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i113 (.D(prev_key0_new_127__N_4659[113]), .SP(clk_c_enable_132), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[113])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i113.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i114 (.D(prev_key0_new_127__N_4659[114]), .SP(clk_c_enable_132), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[114])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i114.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i115 (.D(prev_key0_new_127__N_4659[115]), .SP(clk_c_enable_132), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[115])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i115.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i116 (.D(prev_key0_new_127__N_4659[116]), .SP(clk_c_enable_132), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[116])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i116.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i117 (.D(prev_key0_new_127__N_4659[117]), .SP(clk_c_enable_132), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[117])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i117.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i118 (.D(prev_key0_new_127__N_4659[118]), .SP(clk_c_enable_132), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[118])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i118.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i119 (.D(prev_key0_new_127__N_4659[119]), .SP(clk_c_enable_132), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[119])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i119.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i120 (.D(prev_key0_new_127__N_4659[120]), .SP(clk_c_enable_132), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[120])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i120.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i121 (.D(prev_key0_new_127__N_4659[121]), .SP(clk_c_enable_132), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[121])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i121.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i122 (.D(prev_key0_new_127__N_4659[122]), .SP(clk_c_enable_132), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[122])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i122.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i123 (.D(prev_key0_new_127__N_4659[123]), .SP(clk_c_enable_132), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[123])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i123.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i124 (.D(prev_key0_new_127__N_4659[124]), .SP(clk_c_enable_132), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[124])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i124.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i125 (.D(prev_key0_new_127__N_4659[125]), .SP(clk_c_enable_132), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[125])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i125.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i126 (.D(prev_key0_new_127__N_4659[126]), .SP(clk_c_enable_132), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[126])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i126.GSR = "DISABLED";
    FD1P3IX prev_key0_reg__i127 (.D(prev_key0_new_127__N_4659[127]), .SP(clk_c_enable_132), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key0_reg[127])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key0_reg__i127.GSR = "DISABLED";
    L6MUX21 i25287 (.D0(n30443), .D1(n33404), .SD(\muxed_round_nr[2] ), 
            .Z(n30446));
    LUT4 round_3__I_0_Mux_45_i4_3_lut (.A(\key_mem[4] [45]), .B(\key_mem[5] [45]), 
         .C(maxfan_replicated_net_23), .Z(n4_adj_9195)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_45_i4_3_lut.init = 16'hcaca;
    L6MUX21 i25293 (.D0(n30448), .D1(n30449), .SD(\muxed_round_nr[2] ), 
            .Z(n30452));
    LUT4 round_3__I_0_Mux_45_i2_3_lut (.A(\key_mem[2] [45]), .B(\key_mem[3] [45]), 
         .C(maxfan_replicated_net_23), .Z(n2_adj_9196)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_45_i2_3_lut.init = 16'hcaca;
    L6MUX21 i25294 (.D0(n30450), .D1(n33407), .SD(\muxed_round_nr[2] ), 
            .Z(n30453));
    LUT4 round_3__I_0_Mux_45_i1_3_lut (.A(\key_mem[0] [45]), .B(\key_mem[1] [45]), 
         .C(maxfan_replicated_net_23), .Z(n1_adj_9197)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_45_i1_3_lut.init = 16'hcaca;
    L6MUX21 i25300 (.D0(n30455), .D1(n30456), .SD(\muxed_round_nr[2] ), 
            .Z(n30459));
    LUT4 mux_9_i26_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [25]), 
         .D(key_mem_new[25]), .Z(key_mem_0__127__N_6752[25])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i26_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i27_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [26]), 
         .D(key_mem_new[26]), .Z(key_mem_0__127__N_6752[26])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i27_3_lut_4_lut.init = 16'hf4b0;
    L6MUX21 i25301 (.D0(n30457), .D1(n33408), .SD(\muxed_round_nr[2] ), 
            .Z(n30460));
    L6MUX21 i25307 (.D0(n30462), .D1(n30463), .SD(\muxed_round_nr[2] ), 
            .Z(n30466));
    L6MUX21 i25308 (.D0(n30464), .D1(n33410), .SD(\muxed_round_nr[2] ), 
            .Z(n30467));
    LUT4 mux_9_i28_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [27]), 
         .D(key_mem_new[27]), .Z(key_mem_0__127__N_6752[27])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i28_3_lut_4_lut.init = 16'hf4b0;
    L6MUX21 i25314 (.D0(n30469), .D1(n30470), .SD(\muxed_round_nr[2] ), 
            .Z(n30473));
    LUT4 round_3__I_0_Mux_44_i11_3_lut (.A(\key_mem[12] [44]), .B(\key_mem[13] [44]), 
         .C(maxfan_replicated_net_23), .Z(n11_adj_116)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_44_i11_3_lut.init = 16'hcaca;
    LUT4 i15044_2_lut_4_lut (.A(\key_reg[4] [9]), .B(n4_adj_8349), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[105])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15044_2_lut_4_lut.init = 16'hca00;
    LUT4 round_3__I_0_Mux_44_i9_3_lut (.A(\key_mem[10] [44]), .B(\key_mem[11] [44]), 
         .C(maxfan_replicated_net_23), .Z(n9_adj_9199)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_44_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_44_i8_3_lut (.A(\key_mem[8] [44]), .B(\key_mem[9] [44]), 
         .C(maxfan_replicated_net_23), .Z(n8_adj_9200)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_44_i8_3_lut.init = 16'hcaca;
    L6MUX21 i25315 (.D0(n30471), .D1(n33412), .SD(\muxed_round_nr[2] ), 
            .Z(n30474));
    LUT4 mux_9_i29_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [28]), 
         .D(key_mem_new[28]), .Z(key_mem_0__127__N_6752[28])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i29_3_lut_4_lut.init = 16'hf4b0;
    LUT4 round_3__I_0_Mux_44_i5_3_lut (.A(\key_mem[6] [44]), .B(\key_mem[7] [44]), 
         .C(maxfan_replicated_net_23), .Z(n5_adj_9201)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_44_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_44_i4_3_lut (.A(\key_mem[4] [44]), .B(\key_mem[5] [44]), 
         .C(maxfan_replicated_net_23), .Z(n4_adj_9202)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_44_i4_3_lut.init = 16'hcaca;
    L6MUX21 i25321 (.D0(n30476), .D1(n30477), .SD(\muxed_round_nr[2] ), 
            .Z(n30480));
    L6MUX21 i25322 (.D0(n30478), .D1(n33414), .SD(\muxed_round_nr[2] ), 
            .Z(n30481));
    L6MUX21 i25328 (.D0(n30483), .D1(n30484), .SD(\muxed_round_nr[2] ), 
            .Z(n30487));
    LUT4 round_3__I_0_Mux_44_i2_3_lut (.A(\key_mem[2] [44]), .B(\key_mem[3] [44]), 
         .C(maxfan_replicated_net_23), .Z(n2_adj_9203)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_44_i2_3_lut.init = 16'hcaca;
    L6MUX21 i25329 (.D0(n30485), .D1(n33415), .SD(\muxed_round_nr[2] ), 
            .Z(n30488));
    LUT4 round_3__I_0_Mux_44_i1_3_lut (.A(\key_mem[0] [44]), .B(\key_mem[1] [44]), 
         .C(maxfan_replicated_net_23), .Z(n1_adj_9204)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_44_i1_3_lut.init = 16'hcaca;
    L6MUX21 i25335 (.D0(n30490), .D1(n30491), .SD(\muxed_round_nr[2] ), 
            .Z(n30494));
    LUT4 round_3__I_0_Mux_121_i8_3_lut (.A(\key_mem[8] [121]), .B(\key_mem[9] [121]), 
         .C(n33952), .Z(n8_adj_9205)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_121_i8_3_lut.init = 16'hcaca;
    LUT4 mux_9_i30_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [29]), 
         .D(key_mem_new[29]), .Z(key_mem_0__127__N_6752[29])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i30_3_lut_4_lut.init = 16'hf4b0;
    L6MUX21 i25336 (.D0(n30492), .D1(n33416), .SD(\muxed_round_nr[2] ), 
            .Z(n30495));
    LUT4 mux_9_i31_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [30]), 
         .D(key_mem_new[30]), .Z(key_mem_0__127__N_6752[30])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i31_3_lut_4_lut.init = 16'hf4b0;
    L6MUX21 i25342 (.D0(n30497), .D1(n30498), .SD(\muxed_round_nr[2] ), 
            .Z(n30501));
    LUT4 round_3__I_0_Mux_43_i11_3_lut (.A(\key_mem[12] [43]), .B(\key_mem[13] [43]), 
         .C(maxfan_replicated_net_23), .Z(n11_adj_117)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_43_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_43_i9_3_lut (.A(\key_mem[10] [43]), .B(\key_mem[11] [43]), 
         .C(maxfan_replicated_net_23), .Z(n9_adj_9207)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_43_i9_3_lut.init = 16'hcaca;
    L6MUX21 i25343 (.D0(n30499), .D1(n33417), .SD(\muxed_round_nr[2] ), 
            .Z(n30502));
    LUT4 round_3__I_0_Mux_43_i8_3_lut (.A(\key_mem[8] [43]), .B(\key_mem[9] [43]), 
         .C(maxfan_replicated_net_23), .Z(n8_adj_9208)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_43_i8_3_lut.init = 16'hcaca;
    L6MUX21 i25349 (.D0(n30504), .D1(n30505), .SD(\muxed_round_nr[2] ), 
            .Z(n30508));
    LUT4 round_3__I_0_Mux_43_i5_3_lut (.A(\key_mem[6] [43]), .B(\key_mem[7] [43]), 
         .C(maxfan_replicated_net_23), .Z(n5_adj_9209)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_43_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_43_i4_3_lut (.A(\key_mem[4] [43]), .B(\key_mem[5] [43]), 
         .C(maxfan_replicated_net_23), .Z(n4_adj_9210)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_43_i4_3_lut.init = 16'hcaca;
    L6MUX21 i25350 (.D0(n30506), .D1(n33418), .SD(\muxed_round_nr[2] ), 
            .Z(n30509));
    LUT4 round_3__I_0_Mux_43_i2_3_lut (.A(\key_mem[2] [43]), .B(\key_mem[3] [43]), 
         .C(maxfan_replicated_net_23), .Z(n2_adj_9211)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_43_i2_3_lut.init = 16'hcaca;
    L6MUX21 i25356 (.D0(n30511), .D1(n30512), .SD(\muxed_round_nr[2] ), 
            .Z(n30515));
    LUT4 round_3__I_0_Mux_43_i1_3_lut (.A(\key_mem[0] [43]), .B(\key_mem[1] [43]), 
         .C(maxfan_replicated_net_23), .Z(n1_adj_9212)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_43_i1_3_lut.init = 16'hcaca;
    L6MUX21 i25357 (.D0(n30513), .D1(n33419), .SD(\muxed_round_nr[2] ), 
            .Z(n30516));
    LUT4 round_3__I_0_Mux_25_i2_3_lut (.A(\key_mem[2] [25]), .B(\key_mem[3] [25]), 
         .C(maxfan_replicated_net_23), .Z(n2_adj_9213)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_25_i2_3_lut.init = 16'hcaca;
    L6MUX21 i25363 (.D0(n30518), .D1(n30519), .SD(\muxed_round_nr[2] ), 
            .Z(n30522));
    LUT4 round_3__I_0_Mux_25_i1_3_lut (.A(\key_mem[0] [25]), .B(\key_mem[1] [25]), 
         .C(maxfan_replicated_net_23), .Z(n1_adj_9214)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_25_i1_3_lut.init = 16'hcaca;
    L6MUX21 i25364 (.D0(n30520), .D1(n33420), .SD(\muxed_round_nr[2] ), 
            .Z(n30523));
    L6MUX21 i25370 (.D0(n30525), .D1(n30526), .SD(\muxed_round_nr[2] ), 
            .Z(n30529));
    LUT4 mux_9_i32_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [31]), 
         .D(key_mem_new[31]), .Z(key_mem_0__127__N_6752[31])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i32_3_lut_4_lut.init = 16'hf4b0;
    L6MUX21 i25371 (.D0(n30527), .D1(n33421), .SD(\muxed_round_nr[2] ), 
            .Z(n30530));
    L6MUX21 i25377 (.D0(n30532), .D1(n30533), .SD(\muxed_round_nr[2] ), 
            .Z(n30536));
    LUT4 round_3__I_0_Mux_121_i5_3_lut (.A(\key_mem[6] [121]), .B(\key_mem[7] [121]), 
         .C(n33952), .Z(n5_adj_9215)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_121_i5_3_lut.init = 16'hcaca;
    L6MUX21 i25378 (.D0(n30534), .D1(n33422), .SD(\muxed_round_nr[2] ), 
            .Z(n30537));
    L6MUX21 i25384 (.D0(n30539), .D1(n30540), .SD(\muxed_round_nr[2] ), 
            .Z(n30543));
    L6MUX21 i25385 (.D0(n30541), .D1(n33423), .SD(\muxed_round_nr[2] ), 
            .Z(n30544));
    LUT4 mux_9_i33_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [32]), 
         .D(key_mem_new[32]), .Z(key_mem_0__127__N_6752[32])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i33_3_lut_4_lut.init = 16'hf4b0;
    L6MUX21 i25391 (.D0(n30546), .D1(n30547), .SD(\muxed_round_nr[2] ), 
            .Z(n30550));
    LUT4 mux_9_i34_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [33]), 
         .D(key_mem_new[33]), .Z(key_mem_0__127__N_6752[33])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i34_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i35_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [34]), 
         .D(key_mem_new[34]), .Z(key_mem_0__127__N_6752[34])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i35_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i36_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [35]), 
         .D(key_mem_new[35]), .Z(key_mem_0__127__N_6752[35])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i36_3_lut_4_lut.init = 16'hf4b0;
    L6MUX21 i25392 (.D0(n30548), .D1(n33424), .SD(\muxed_round_nr[2] ), 
            .Z(n30551));
    LUT4 mux_9_i37_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [36]), 
         .D(key_mem_new[36]), .Z(key_mem_0__127__N_6752[36])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i37_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i38_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [37]), 
         .D(key_mem_new[37]), .Z(key_mem_0__127__N_6752[37])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i38_3_lut_4_lut.init = 16'hf4b0;
    L6MUX21 i25398 (.D0(n30553), .D1(n30554), .SD(\muxed_round_nr[2] ), 
            .Z(n30557));
    LUT4 round_3__I_0_Mux_121_i4_3_lut (.A(\key_mem[4] [121]), .B(\key_mem[5] [121]), 
         .C(n33952), .Z(n4_adj_9216)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_121_i4_3_lut.init = 16'hcaca;
    L6MUX21 i25399 (.D0(n30555), .D1(n33425), .SD(\muxed_round_nr[2] ), 
            .Z(n30558));
    LUT4 mux_9_i39_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [38]), 
         .D(key_mem_new[38]), .Z(key_mem_0__127__N_6752[38])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i39_3_lut_4_lut.init = 16'hf4b0;
    L6MUX21 i25405 (.D0(n30560), .D1(n30561), .SD(\muxed_round_nr[2] ), 
            .Z(n30564));
    LUT4 mux_9_i66_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [65]), 
         .D(key_mem_new[65]), .Z(key_mem_0__127__N_6752[65])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i66_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i67_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [66]), 
         .D(key_mem_new[66]), .Z(key_mem_0__127__N_6752[66])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i67_3_lut_4_lut.init = 16'hf4b0;
    L6MUX21 i25406 (.D0(n30562), .D1(n33426), .SD(\muxed_round_nr[2] ), 
            .Z(n30565));
    LUT4 mux_9_i68_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [67]), 
         .D(key_mem_new[67]), .Z(key_mem_0__127__N_6752[67])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i68_3_lut_4_lut.init = 16'hf4b0;
    L6MUX21 i25412 (.D0(n30567), .D1(n30568), .SD(\muxed_round_nr[2] ), 
            .Z(n30571));
    FD1P3AX rcon_reg_i0_i2 (.D(rcon_new[2]), .SP(rcon_we), .CK(clk_c), 
            .Q(rcon_reg[2])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam rcon_reg_i0_i2.GSR = "ENABLED";
    FD1P3AX rcon_reg_i0_i3 (.D(rcon_new[3]), .SP(rcon_we), .CK(clk_c), 
            .Q(rcon_reg[3])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam rcon_reg_i0_i3.GSR = "ENABLED";
    LUT4 round_3__I_0_Mux_104_i4_3_lut (.A(\key_mem[4] [104]), .B(\key_mem[5] [104]), 
         .C(n33952), .Z(n4_adj_9217)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_104_i4_3_lut.init = 16'hcaca;
    LUT4 mux_9_i69_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [68]), 
         .D(key_mem_new[68]), .Z(key_mem_0__127__N_6752[68])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i69_3_lut_4_lut.init = 16'hf4b0;
    FD1P3AX rcon_reg_i0_i7 (.D(rcon_new[7]), .SP(rcon_we), .CK(clk_c), 
            .Q(\rcon_logic.tmp_rcon [0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam rcon_reg_i0_i7.GSR = "ENABLED";
    L6MUX21 i25413 (.D0(n30569), .D1(n33427), .SD(\muxed_round_nr[2] ), 
            .Z(n30572));
    LUT4 mux_9_i70_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [69]), 
         .D(key_mem_new[69]), .Z(key_mem_0__127__N_6752[69])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i70_3_lut_4_lut.init = 16'hf4b0;
    L6MUX21 i25419 (.D0(n30574), .D1(n30575), .SD(\muxed_round_nr[2] ), 
            .Z(n30578));
    LUT4 mux_9_i71_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [70]), 
         .D(key_mem_new[70]), .Z(key_mem_0__127__N_6752[70])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i71_3_lut_4_lut.init = 16'hf4b0;
    L6MUX21 i25420 (.D0(n30576), .D1(n33428), .SD(\muxed_round_nr[2] ), 
            .Z(n30579));
    LUT4 mux_9_i72_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [71]), 
         .D(key_mem_new[71]), .Z(key_mem_0__127__N_6752[71])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i72_3_lut_4_lut.init = 16'hf4b0;
    LUT4 round_3__I_0_Mux_104_i2_3_lut (.A(\key_mem[2] [104]), .B(\key_mem[3] [104]), 
         .C(n33952), .Z(n2_adj_9218)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_104_i2_3_lut.init = 16'hcaca;
    LUT4 mux_9_i73_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [72]), 
         .D(key_mem_new[72]), .Z(key_mem_0__127__N_6752[72])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i73_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i74_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [73]), 
         .D(key_mem_new[73]), .Z(key_mem_0__127__N_6752[73])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i74_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i75_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [74]), 
         .D(key_mem_new[74]), .Z(key_mem_0__127__N_6752[74])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i75_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i76_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [75]), 
         .D(key_mem_new[75]), .Z(key_mem_0__127__N_6752[75])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i76_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i77_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [76]), 
         .D(key_mem_new[76]), .Z(key_mem_0__127__N_6752[76])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i77_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i78_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [77]), 
         .D(key_mem_new[77]), .Z(key_mem_0__127__N_6752[77])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i78_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i79_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [78]), 
         .D(key_mem_new[78]), .Z(key_mem_0__127__N_6752[78])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i79_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i80_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [79]), 
         .D(key_mem_new[79]), .Z(key_mem_0__127__N_6752[79])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i80_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i81_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [80]), 
         .D(key_mem_new[80]), .Z(key_mem_0__127__N_6752[80])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i81_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i82_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [81]), 
         .D(key_mem_new[81]), .Z(key_mem_0__127__N_6752[81])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i82_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i83_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [82]), 
         .D(key_mem_new[82]), .Z(key_mem_0__127__N_6752[82])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i83_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i84_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [83]), 
         .D(key_mem_new[83]), .Z(key_mem_0__127__N_6752[83])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i84_3_lut_4_lut.init = 16'hf4b0;
    LUT4 round_3__I_0_Mux_104_i1_3_lut (.A(\key_mem[0] [104]), .B(\key_mem[1] [104]), 
         .C(n33952), .Z(n1_adj_9219)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_104_i1_3_lut.init = 16'hcaca;
    LUT4 mux_9_i85_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [84]), 
         .D(key_mem_new[84]), .Z(key_mem_0__127__N_6752[84])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i85_3_lut_4_lut.init = 16'hf4b0;
    L6MUX21 i25426 (.D0(n30581), .D1(n30582), .SD(\muxed_round_nr[2] ), 
            .Z(n30585));
    LUT4 mux_9_i86_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [85]), 
         .D(key_mem_new[85]), .Z(key_mem_0__127__N_6752[85])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i86_3_lut_4_lut.init = 16'hf4b0;
    L6MUX21 i25427 (.D0(n30583), .D1(n33429), .SD(\muxed_round_nr[2] ), 
            .Z(n30586));
    LUT4 mux_9_i87_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [86]), 
         .D(key_mem_new[86]), .Z(key_mem_0__127__N_6752[86])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i87_3_lut_4_lut.init = 16'hf4b0;
    L6MUX21 i25433 (.D0(n30588), .D1(n30589), .SD(\muxed_round_nr[2] ), 
            .Z(n30592));
    LUT4 mux_9_i88_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [87]), 
         .D(key_mem_new[87]), .Z(key_mem_0__127__N_6752[87])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i88_3_lut_4_lut.init = 16'hf4b0;
    L6MUX21 i25434 (.D0(n30590), .D1(n33430), .SD(\muxed_round_nr[2] ), 
            .Z(n30593));
    LUT4 mux_9_i89_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [88]), 
         .D(key_mem_new[88]), .Z(key_mem_0__127__N_6752[88])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i89_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i90_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [89]), 
         .D(key_mem_new[89]), .Z(key_mem_0__127__N_6752[89])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i90_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i91_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [90]), 
         .D(key_mem_new[90]), .Z(key_mem_0__127__N_6752[90])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i91_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i92_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [91]), 
         .D(key_mem_new[91]), .Z(key_mem_0__127__N_6752[91])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i92_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i93_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [92]), 
         .D(key_mem_new[92]), .Z(key_mem_0__127__N_6752[92])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i93_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i94_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [93]), 
         .D(key_mem_new[93]), .Z(key_mem_0__127__N_6752[93])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i94_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i95_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [94]), 
         .D(key_mem_new[94]), .Z(key_mem_0__127__N_6752[94])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i95_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i96_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [95]), 
         .D(key_mem_new[95]), .Z(key_mem_0__127__N_6752[95])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i96_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i97_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [96]), 
         .D(key_mem_new[96]), .Z(key_mem_0__127__N_6752[96])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i97_3_lut_4_lut.init = 16'hf4b0;
    L6MUX21 i25440 (.D0(n30595), .D1(n30596), .SD(\muxed_round_nr[2] ), 
            .Z(n30599));
    LUT4 mux_9_i98_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [97]), 
         .D(key_mem_new[97]), .Z(key_mem_0__127__N_6752[97])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i98_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i99_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [98]), 
         .D(key_mem_new[98]), .Z(key_mem_0__127__N_6752[98])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i99_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i100_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [99]), 
         .D(key_mem_new[99]), .Z(key_mem_0__127__N_6752[99])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i100_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i101_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [100]), 
         .D(key_mem_new[100]), .Z(key_mem_0__127__N_6752[100])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i101_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i102_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [101]), 
         .D(key_mem_new[101]), .Z(key_mem_0__127__N_6752[101])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i102_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i103_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [102]), 
         .D(key_mem_new[102]), .Z(key_mem_0__127__N_6752[102])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i103_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i104_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [103]), 
         .D(key_mem_new[103]), .Z(key_mem_0__127__N_6752[103])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i104_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i105_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [104]), 
         .D(key_mem_new[104]), .Z(key_mem_0__127__N_6752[104])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i105_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i106_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [105]), 
         .D(key_mem_new[105]), .Z(key_mem_0__127__N_6752[105])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i106_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i107_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [106]), 
         .D(key_mem_new[106]), .Z(key_mem_0__127__N_6752[106])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i107_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i108_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [107]), 
         .D(key_mem_new[107]), .Z(key_mem_0__127__N_6752[107])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i108_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i109_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [108]), 
         .D(key_mem_new[108]), .Z(key_mem_0__127__N_6752[108])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i109_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i110_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [109]), 
         .D(key_mem_new[109]), .Z(key_mem_0__127__N_6752[109])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i110_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i111_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [110]), 
         .D(key_mem_new[110]), .Z(key_mem_0__127__N_6752[110])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i111_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i112_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [111]), 
         .D(key_mem_new[111]), .Z(key_mem_0__127__N_6752[111])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i112_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i113_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [112]), 
         .D(key_mem_new[112]), .Z(key_mem_0__127__N_6752[112])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i113_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i114_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [113]), 
         .D(key_mem_new[113]), .Z(key_mem_0__127__N_6752[113])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i114_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i115_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [114]), 
         .D(key_mem_new[114]), .Z(key_mem_0__127__N_6752[114])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i115_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i116_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [115]), 
         .D(key_mem_new[115]), .Z(key_mem_0__127__N_6752[115])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i116_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i117_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [116]), 
         .D(key_mem_new[116]), .Z(key_mem_0__127__N_6752[116])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i117_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i118_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [117]), 
         .D(key_mem_new[117]), .Z(key_mem_0__127__N_6752[117])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i118_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i119_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [118]), 
         .D(key_mem_new[118]), .Z(key_mem_0__127__N_6752[118])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i119_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i120_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [119]), 
         .D(key_mem_new[119]), .Z(key_mem_0__127__N_6752[119])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i120_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i121_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [120]), 
         .D(key_mem_new[120]), .Z(key_mem_0__127__N_6752[120])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i121_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i122_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [121]), 
         .D(key_mem_new[121]), .Z(key_mem_0__127__N_6752[121])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i122_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i123_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [122]), 
         .D(key_mem_new[122]), .Z(key_mem_0__127__N_6752[122])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i123_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i124_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [123]), 
         .D(key_mem_new[123]), .Z(key_mem_0__127__N_6752[123])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i124_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i125_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [124]), 
         .D(key_mem_new[124]), .Z(key_mem_0__127__N_6752[124])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i125_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i126_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [125]), 
         .D(key_mem_new[125]), .Z(key_mem_0__127__N_6752[125])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i126_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i127_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [126]), 
         .D(key_mem_new[126]), .Z(key_mem_0__127__N_6752[126])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i127_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i128_3_lut_4_lut (.A(n33912), .B(n33911), .C(\key_mem[14] [127]), 
         .D(key_mem_new[127]), .Z(key_mem_0__127__N_6752[127])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_9_i128_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_21_i1_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [0]), 
         .D(key_mem_new[0]), .Z(key_mem_0__127__N_5216[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i2_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [1]), 
         .D(key_mem_new[1]), .Z(key_mem_0__127__N_5216[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i3_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [2]), 
         .D(key_mem_new[2]), .Z(key_mem_0__127__N_5216[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i4_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [3]), 
         .D(key_mem_new[3]), .Z(key_mem_0__127__N_5216[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i5_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [4]), 
         .D(key_mem_new[4]), .Z(key_mem_0__127__N_5216[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i6_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [5]), 
         .D(key_mem_new[5]), .Z(key_mem_0__127__N_5216[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i7_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [6]), 
         .D(key_mem_new[6]), .Z(key_mem_0__127__N_5216[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i8_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [7]), 
         .D(key_mem_new[7]), .Z(key_mem_0__127__N_5216[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i9_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [8]), 
         .D(key_mem_new[8]), .Z(key_mem_0__127__N_5216[8])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i9_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i10_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [9]), 
         .D(key_mem_new[9]), .Z(key_mem_0__127__N_5216[9])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i10_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i11_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [10]), 
         .D(key_mem_new[10]), .Z(key_mem_0__127__N_5216[10])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i11_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i12_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [11]), 
         .D(key_mem_new[11]), .Z(key_mem_0__127__N_5216[11])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i12_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i13_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [12]), 
         .D(key_mem_new[12]), .Z(key_mem_0__127__N_5216[12])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i13_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i14_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [13]), 
         .D(key_mem_new[13]), .Z(key_mem_0__127__N_5216[13])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i14_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i15_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [14]), 
         .D(key_mem_new[14]), .Z(key_mem_0__127__N_5216[14])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i15_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i16_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [15]), 
         .D(key_mem_new[15]), .Z(key_mem_0__127__N_5216[15])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i16_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i17_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [16]), 
         .D(key_mem_new[16]), .Z(key_mem_0__127__N_5216[16])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i17_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i18_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [17]), 
         .D(key_mem_new[17]), .Z(key_mem_0__127__N_5216[17])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i18_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i19_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [18]), 
         .D(key_mem_new[18]), .Z(key_mem_0__127__N_5216[18])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i19_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i20_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [19]), 
         .D(key_mem_new[19]), .Z(key_mem_0__127__N_5216[19])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i20_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i21_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [20]), 
         .D(key_mem_new[20]), .Z(key_mem_0__127__N_5216[20])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i21_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i22_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [21]), 
         .D(key_mem_new[21]), .Z(key_mem_0__127__N_5216[21])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i22_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i23_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [22]), 
         .D(key_mem_new[22]), .Z(key_mem_0__127__N_5216[22])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i23_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i24_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [23]), 
         .D(key_mem_new[23]), .Z(key_mem_0__127__N_5216[23])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i24_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i25_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [24]), 
         .D(key_mem_new[24]), .Z(key_mem_0__127__N_5216[24])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i25_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i26_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [25]), 
         .D(key_mem_new[25]), .Z(key_mem_0__127__N_5216[25])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i26_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i27_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [26]), 
         .D(key_mem_new[26]), .Z(key_mem_0__127__N_5216[26])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i27_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i28_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [27]), 
         .D(key_mem_new[27]), .Z(key_mem_0__127__N_5216[27])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i28_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i29_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [28]), 
         .D(key_mem_new[28]), .Z(key_mem_0__127__N_5216[28])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i29_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i30_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [29]), 
         .D(key_mem_new[29]), .Z(key_mem_0__127__N_5216[29])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i30_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i31_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [30]), 
         .D(key_mem_new[30]), .Z(key_mem_0__127__N_5216[30])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i31_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i32_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [31]), 
         .D(key_mem_new[31]), .Z(key_mem_0__127__N_5216[31])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i32_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i33_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [32]), 
         .D(key_mem_new[32]), .Z(key_mem_0__127__N_5216[32])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i33_3_lut_4_lut.init = 16'hf1e0;
    LUT4 round_3__I_0_Mux_121_i2_3_lut (.A(\key_mem[2] [121]), .B(\key_mem[3] [121]), 
         .C(n33952), .Z(n2_adj_9220)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_121_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_121_i1_3_lut (.A(\key_mem[0] [121]), .B(\key_mem[1] [121]), 
         .C(n33952), .Z(n1_adj_9221)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_121_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_120_i11_3_lut (.A(\key_mem[12] [120]), .B(\key_mem[13] [120]), 
         .C(n33952), .Z(n11_adj_118)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_120_i11_3_lut.init = 16'hcaca;
    LUT4 mux_21_i34_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [33]), 
         .D(key_mem_new[33]), .Z(key_mem_0__127__N_5216[33])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i34_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15043_2_lut_4_lut (.A(\key_reg[4] [8]), .B(n4_adj_8343), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[104])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15043_2_lut_4_lut.init = 16'hca00;
    LUT4 round_3__I_0_Mux_120_i9_3_lut (.A(\key_mem[10] [120]), .B(\key_mem[11] [120]), 
         .C(n33952), .Z(n9_adj_9223)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_120_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_120_i8_3_lut (.A(\key_mem[8] [120]), .B(\key_mem[9] [120]), 
         .C(n33952), .Z(n8_adj_9224)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_120_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_120_i5_3_lut (.A(\key_mem[6] [120]), .B(\key_mem[7] [120]), 
         .C(n33952), .Z(n5_adj_9225)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_120_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_120_i4_3_lut (.A(\key_mem[4] [120]), .B(\key_mem[5] [120]), 
         .C(n33952), .Z(n4_adj_9226)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_120_i4_3_lut.init = 16'hcaca;
    LUT4 mux_21_i35_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [34]), 
         .D(key_mem_new[34]), .Z(key_mem_0__127__N_5216[34])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i35_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i36_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [35]), 
         .D(key_mem_new[35]), .Z(key_mem_0__127__N_5216[35])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i36_3_lut_4_lut.init = 16'hf1e0;
    LUT4 round_3__I_0_Mux_120_i2_3_lut (.A(\key_mem[2] [120]), .B(\key_mem[3] [120]), 
         .C(n33952), .Z(n2_adj_9227)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_120_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_120_i1_3_lut (.A(\key_mem[0] [120]), .B(\key_mem[1] [120]), 
         .C(n33952), .Z(n1_adj_9228)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_120_i1_3_lut.init = 16'hcaca;
    LUT4 mux_21_i37_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [36]), 
         .D(key_mem_new[36]), .Z(key_mem_0__127__N_5216[36])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i37_3_lut_4_lut.init = 16'hf1e0;
    LUT4 round_3__I_0_Mux_119_i11_3_lut (.A(\key_mem[12] [119]), .B(\key_mem[13] [119]), 
         .C(n33952), .Z(n11_adj_119)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_119_i11_3_lut.init = 16'hcaca;
    LUT4 mux_21_i38_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [37]), 
         .D(key_mem_new[37]), .Z(key_mem_0__127__N_5216[37])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i38_3_lut_4_lut.init = 16'hf1e0;
    LUT4 round_3__I_0_Mux_119_i9_3_lut (.A(\key_mem[10] [119]), .B(\key_mem[11] [119]), 
         .C(n33952), .Z(n9_adj_9230)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_119_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_119_i8_3_lut (.A(\key_mem[8] [119]), .B(\key_mem[9] [119]), 
         .C(n33952), .Z(n8_adj_9231)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_119_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_119_i5_3_lut (.A(\key_mem[6] [119]), .B(\key_mem[7] [119]), 
         .C(n33952), .Z(n5_adj_9232)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_119_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_119_i4_3_lut (.A(\key_mem[4] [119]), .B(\key_mem[5] [119]), 
         .C(n33952), .Z(n4_adj_9233)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_119_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_119_i2_3_lut (.A(\key_mem[2] [119]), .B(\key_mem[3] [119]), 
         .C(n33952), .Z(n2_adj_9234)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_119_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_119_i1_3_lut (.A(\key_mem[0] [119]), .B(\key_mem[1] [119]), 
         .C(n33952), .Z(n1_adj_9235)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_119_i1_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_118_i11_3_lut (.A(\key_mem[12] [118]), .B(\key_mem[13] [118]), 
         .C(n33952), .Z(n11_adj_120)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_118_i11_3_lut.init = 16'hcaca;
    LUT4 i15042_2_lut_4_lut (.A(\key_reg[4] [7]), .B(n4_adj_8339), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[103])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15042_2_lut_4_lut.init = 16'hca00;
    LUT4 round_3__I_0_Mux_118_i9_3_lut (.A(\key_mem[10] [118]), .B(\key_mem[11] [118]), 
         .C(n33952), .Z(n9_adj_9237)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_118_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_118_i8_3_lut (.A(\key_mem[8] [118]), .B(\key_mem[9] [118]), 
         .C(n33952), .Z(n8_adj_9238)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_118_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_118_i5_3_lut (.A(\key_mem[6] [118]), .B(\key_mem[7] [118]), 
         .C(n33952), .Z(n5_adj_9239)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_118_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_118_i4_3_lut (.A(\key_mem[4] [118]), .B(\key_mem[5] [118]), 
         .C(n33952), .Z(n4_adj_9240)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_118_i4_3_lut.init = 16'hcaca;
    LUT4 mux_21_i39_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [38]), 
         .D(key_mem_new[38]), .Z(key_mem_0__127__N_5216[38])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i39_3_lut_4_lut.init = 16'hf1e0;
    LUT4 round_3__I_0_Mux_118_i2_3_lut (.A(\key_mem[2] [118]), .B(\key_mem[3] [118]), 
         .C(n33952), .Z(n2_adj_9241)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_118_i2_3_lut.init = 16'hcaca;
    LUT4 mux_21_i40_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [39]), 
         .D(key_mem_new[39]), .Z(key_mem_0__127__N_5216[39])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i40_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i41_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [40]), 
         .D(key_mem_new[40]), .Z(key_mem_0__127__N_5216[40])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i41_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i42_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [41]), 
         .D(key_mem_new[41]), .Z(key_mem_0__127__N_5216[41])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i42_3_lut_4_lut.init = 16'hf1e0;
    LUT4 round_3__I_0_Mux_118_i1_3_lut (.A(\key_mem[0] [118]), .B(\key_mem[1] [118]), 
         .C(n33952), .Z(n1_adj_9242)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_118_i1_3_lut.init = 16'hcaca;
    LUT4 mux_21_i43_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [42]), 
         .D(key_mem_new[42]), .Z(key_mem_0__127__N_5216[42])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i43_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i44_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [43]), 
         .D(key_mem_new[43]), .Z(key_mem_0__127__N_5216[43])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i44_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i45_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [44]), 
         .D(key_mem_new[44]), .Z(key_mem_0__127__N_5216[44])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i45_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i46_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [45]), 
         .D(key_mem_new[45]), .Z(key_mem_0__127__N_5216[45])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i46_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i47_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [46]), 
         .D(key_mem_new[46]), .Z(key_mem_0__127__N_5216[46])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i47_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i48_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [47]), 
         .D(key_mem_new[47]), .Z(key_mem_0__127__N_5216[47])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i48_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i49_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [48]), 
         .D(key_mem_new[48]), .Z(key_mem_0__127__N_5216[48])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i49_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i50_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [49]), 
         .D(key_mem_new[49]), .Z(key_mem_0__127__N_5216[49])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i50_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i51_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [50]), 
         .D(key_mem_new[50]), .Z(key_mem_0__127__N_5216[50])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i51_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i52_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [51]), 
         .D(key_mem_new[51]), .Z(key_mem_0__127__N_5216[51])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i52_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i53_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [52]), 
         .D(key_mem_new[52]), .Z(key_mem_0__127__N_5216[52])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i53_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i54_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [53]), 
         .D(key_mem_new[53]), .Z(key_mem_0__127__N_5216[53])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i54_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i55_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [54]), 
         .D(key_mem_new[54]), .Z(key_mem_0__127__N_5216[54])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i55_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i56_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [55]), 
         .D(key_mem_new[55]), .Z(key_mem_0__127__N_5216[55])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i56_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i57_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [56]), 
         .D(key_mem_new[56]), .Z(key_mem_0__127__N_5216[56])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i57_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i58_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [57]), 
         .D(key_mem_new[57]), .Z(key_mem_0__127__N_5216[57])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i58_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i59_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [58]), 
         .D(key_mem_new[58]), .Z(key_mem_0__127__N_5216[58])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i59_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i60_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [59]), 
         .D(key_mem_new[59]), .Z(key_mem_0__127__N_5216[59])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i60_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i61_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [60]), 
         .D(key_mem_new[60]), .Z(key_mem_0__127__N_5216[60])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i61_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i62_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [61]), 
         .D(key_mem_new[61]), .Z(key_mem_0__127__N_5216[61])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i62_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i63_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [62]), 
         .D(key_mem_new[62]), .Z(key_mem_0__127__N_5216[62])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i63_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i64_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [63]), 
         .D(key_mem_new[63]), .Z(key_mem_0__127__N_5216[63])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i64_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i65_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [64]), 
         .D(key_mem_new[64]), .Z(key_mem_0__127__N_5216[64])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i65_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i66_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [65]), 
         .D(key_mem_new[65]), .Z(key_mem_0__127__N_5216[65])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i66_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i67_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [66]), 
         .D(key_mem_new[66]), .Z(key_mem_0__127__N_5216[66])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i67_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i68_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [67]), 
         .D(key_mem_new[67]), .Z(key_mem_0__127__N_5216[67])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i68_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i69_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [68]), 
         .D(key_mem_new[68]), .Z(key_mem_0__127__N_5216[68])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i69_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i70_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [69]), 
         .D(key_mem_new[69]), .Z(key_mem_0__127__N_5216[69])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i70_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i71_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [70]), 
         .D(key_mem_new[70]), .Z(key_mem_0__127__N_5216[70])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i71_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i72_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [71]), 
         .D(key_mem_new[71]), .Z(key_mem_0__127__N_5216[71])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i72_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i73_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [72]), 
         .D(key_mem_new[72]), .Z(key_mem_0__127__N_5216[72])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i73_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i74_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [73]), 
         .D(key_mem_new[73]), .Z(key_mem_0__127__N_5216[73])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i74_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i75_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [74]), 
         .D(key_mem_new[74]), .Z(key_mem_0__127__N_5216[74])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i75_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i76_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [75]), 
         .D(key_mem_new[75]), .Z(key_mem_0__127__N_5216[75])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i76_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i77_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [76]), 
         .D(key_mem_new[76]), .Z(key_mem_0__127__N_5216[76])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i77_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i78_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [77]), 
         .D(key_mem_new[77]), .Z(key_mem_0__127__N_5216[77])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i78_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i79_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [78]), 
         .D(key_mem_new[78]), .Z(key_mem_0__127__N_5216[78])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i79_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i80_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [79]), 
         .D(key_mem_new[79]), .Z(key_mem_0__127__N_5216[79])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i80_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i81_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [80]), 
         .D(key_mem_new[80]), .Z(key_mem_0__127__N_5216[80])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i81_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i82_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [81]), 
         .D(key_mem_new[81]), .Z(key_mem_0__127__N_5216[81])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i82_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i83_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [82]), 
         .D(key_mem_new[82]), .Z(key_mem_0__127__N_5216[82])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i83_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i84_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [83]), 
         .D(key_mem_new[83]), .Z(key_mem_0__127__N_5216[83])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i84_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i85_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [84]), 
         .D(key_mem_new[84]), .Z(key_mem_0__127__N_5216[84])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i85_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i86_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [85]), 
         .D(key_mem_new[85]), .Z(key_mem_0__127__N_5216[85])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i86_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i87_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [86]), 
         .D(key_mem_new[86]), .Z(key_mem_0__127__N_5216[86])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i87_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i88_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [87]), 
         .D(key_mem_new[87]), .Z(key_mem_0__127__N_5216[87])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i88_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i89_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [88]), 
         .D(key_mem_new[88]), .Z(key_mem_0__127__N_5216[88])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i89_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i90_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [89]), 
         .D(key_mem_new[89]), .Z(key_mem_0__127__N_5216[89])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i90_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i91_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [90]), 
         .D(key_mem_new[90]), .Z(key_mem_0__127__N_5216[90])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i91_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i92_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [91]), 
         .D(key_mem_new[91]), .Z(key_mem_0__127__N_5216[91])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i92_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i93_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [92]), 
         .D(key_mem_new[92]), .Z(key_mem_0__127__N_5216[92])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i93_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i94_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [93]), 
         .D(key_mem_new[93]), .Z(key_mem_0__127__N_5216[93])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i94_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i95_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [94]), 
         .D(key_mem_new[94]), .Z(key_mem_0__127__N_5216[94])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i95_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i96_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [95]), 
         .D(key_mem_new[95]), .Z(key_mem_0__127__N_5216[95])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i96_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i97_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [96]), 
         .D(key_mem_new[96]), .Z(key_mem_0__127__N_5216[96])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i97_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i98_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [97]), 
         .D(key_mem_new[97]), .Z(key_mem_0__127__N_5216[97])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i98_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i99_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [98]), 
         .D(key_mem_new[98]), .Z(key_mem_0__127__N_5216[98])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i99_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i100_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [99]), 
         .D(key_mem_new[99]), .Z(key_mem_0__127__N_5216[99])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i100_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i101_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [100]), 
         .D(key_mem_new[100]), .Z(key_mem_0__127__N_5216[100])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i101_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i102_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [101]), 
         .D(key_mem_new[101]), .Z(key_mem_0__127__N_5216[101])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i102_3_lut_4_lut.init = 16'hf1e0;
    LUT4 round_3__I_0_Mux_117_i11_3_lut (.A(\key_mem[12] [117]), .B(\key_mem[13] [117]), 
         .C(n33952), .Z(n11_adj_121)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_117_i11_3_lut.init = 16'hcaca;
    LUT4 mux_21_i103_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [102]), 
         .D(key_mem_new[102]), .Z(key_mem_0__127__N_5216[102])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i103_3_lut_4_lut.init = 16'hf1e0;
    LUT4 round_3__I_0_Mux_117_i9_3_lut (.A(\key_mem[10] [117]), .B(\key_mem[11] [117]), 
         .C(n33952), .Z(n9_adj_9244)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_117_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_117_i8_3_lut (.A(\key_mem[8] [117]), .B(\key_mem[9] [117]), 
         .C(n33952), .Z(n8_adj_9245)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_117_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_117_i5_3_lut (.A(\key_mem[6] [117]), .B(\key_mem[7] [117]), 
         .C(n33952), .Z(n5_adj_9246)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_117_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_117_i4_3_lut (.A(\key_mem[4] [117]), .B(\key_mem[5] [117]), 
         .C(n33952), .Z(n4_adj_9247)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_117_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_117_i2_3_lut (.A(\key_mem[2] [117]), .B(\key_mem[3] [117]), 
         .C(n33952), .Z(n2_adj_9248)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_117_i2_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_117_i1_3_lut (.A(\key_mem[0] [117]), .B(\key_mem[1] [117]), 
         .C(n33952), .Z(n1_adj_9249)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_117_i1_3_lut.init = 16'hcaca;
    LUT4 mux_21_i104_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [103]), 
         .D(key_mem_new[103]), .Z(key_mem_0__127__N_5216[103])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i104_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i105_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [104]), 
         .D(key_mem_new[104]), .Z(key_mem_0__127__N_5216[104])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i105_3_lut_4_lut.init = 16'hf1e0;
    LUT4 round_3__I_0_Mux_116_i11_3_lut (.A(\key_mem[12] [116]), .B(\key_mem[13] [116]), 
         .C(n33952), .Z(n11_adj_122)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_116_i11_3_lut.init = 16'hcaca;
    LUT4 i15041_2_lut_4_lut (.A(\key_reg[4] [6]), .B(n4_adj_8337), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[102])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15041_2_lut_4_lut.init = 16'hca00;
    LUT4 round_3__I_0_Mux_116_i9_3_lut (.A(\key_mem[10] [116]), .B(\key_mem[11] [116]), 
         .C(n33952), .Z(n9_adj_9251)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_116_i9_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_116_i8_3_lut (.A(\key_mem[8] [116]), .B(\key_mem[9] [116]), 
         .C(n33952), .Z(n8_adj_9252)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_116_i8_3_lut.init = 16'hcaca;
    LUT4 mux_21_i106_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [105]), 
         .D(key_mem_new[105]), .Z(key_mem_0__127__N_5216[105])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i106_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i107_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [106]), 
         .D(key_mem_new[106]), .Z(key_mem_0__127__N_5216[106])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i107_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i108_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [107]), 
         .D(key_mem_new[107]), .Z(key_mem_0__127__N_5216[107])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i108_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i109_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [108]), 
         .D(key_mem_new[108]), .Z(key_mem_0__127__N_5216[108])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i109_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i110_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [109]), 
         .D(key_mem_new[109]), .Z(key_mem_0__127__N_5216[109])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i110_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i111_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [110]), 
         .D(key_mem_new[110]), .Z(key_mem_0__127__N_5216[110])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i111_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i112_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [111]), 
         .D(key_mem_new[111]), .Z(key_mem_0__127__N_5216[111])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i112_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i113_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [112]), 
         .D(key_mem_new[112]), .Z(key_mem_0__127__N_5216[112])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i113_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i114_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [113]), 
         .D(key_mem_new[113]), .Z(key_mem_0__127__N_5216[113])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i114_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i115_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [114]), 
         .D(key_mem_new[114]), .Z(key_mem_0__127__N_5216[114])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i115_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i116_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [115]), 
         .D(key_mem_new[115]), .Z(key_mem_0__127__N_5216[115])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i116_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i117_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [116]), 
         .D(key_mem_new[116]), .Z(key_mem_0__127__N_5216[116])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i117_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i118_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [117]), 
         .D(key_mem_new[117]), .Z(key_mem_0__127__N_5216[117])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i118_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i119_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [118]), 
         .D(key_mem_new[118]), .Z(key_mem_0__127__N_5216[118])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i119_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i120_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [119]), 
         .D(key_mem_new[119]), .Z(key_mem_0__127__N_5216[119])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i120_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i121_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [120]), 
         .D(key_mem_new[120]), .Z(key_mem_0__127__N_5216[120])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i121_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i122_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [121]), 
         .D(key_mem_new[121]), .Z(key_mem_0__127__N_5216[121])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i122_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i123_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [122]), 
         .D(key_mem_new[122]), .Z(key_mem_0__127__N_5216[122])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i123_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i124_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [123]), 
         .D(key_mem_new[123]), .Z(key_mem_0__127__N_5216[123])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i124_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i125_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [124]), 
         .D(key_mem_new[124]), .Z(key_mem_0__127__N_5216[124])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i125_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i126_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [125]), 
         .D(key_mem_new[125]), .Z(key_mem_0__127__N_5216[125])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i126_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i127_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [126]), 
         .D(key_mem_new[126]), .Z(key_mem_0__127__N_5216[126])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i127_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i128_3_lut_4_lut (.A(n33912), .B(n33944), .C(\key_mem[2] [127]), 
         .D(key_mem_new[127]), .Z(key_mem_0__127__N_5216[127])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_21_i128_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_20_i1_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [0]), 
         .D(key_mem_new[0]), .Z(key_mem_0__127__N_5344[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i1_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i2_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [1]), 
         .D(key_mem_new[1]), .Z(key_mem_0__127__N_5344[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i2_3_lut_4_lut.init = 16'hf2d0;
    FD1P3AX key_mem_14___i2 (.D(key_mem_0__127__N_6752[1]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [1])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i2.GSR = "ENABLED";
    FD1P3AX key_mem_14___i3 (.D(key_mem_0__127__N_6752[2]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [2])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i3.GSR = "ENABLED";
    FD1P3AX key_mem_14___i4 (.D(key_mem_0__127__N_6752[3]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [3])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i4.GSR = "ENABLED";
    FD1P3AX key_mem_14___i5 (.D(key_mem_0__127__N_6752[4]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [4])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i5.GSR = "ENABLED";
    FD1P3AX key_mem_14___i6 (.D(key_mem_0__127__N_6752[5]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [5])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i6.GSR = "ENABLED";
    FD1P3AX key_mem_14___i7 (.D(key_mem_0__127__N_6752[6]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [6])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i7.GSR = "ENABLED";
    FD1P3AX key_mem_14___i8 (.D(key_mem_0__127__N_6752[7]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [7])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i8.GSR = "ENABLED";
    FD1P3AX key_mem_14___i9 (.D(key_mem_0__127__N_6752[8]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [8])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i9.GSR = "ENABLED";
    FD1P3AX key_mem_14___i10 (.D(key_mem_0__127__N_6752[9]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [9])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i10.GSR = "ENABLED";
    FD1P3AX key_mem_14___i11 (.D(key_mem_0__127__N_6752[10]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [10])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i11.GSR = "ENABLED";
    FD1P3AX key_mem_14___i12 (.D(key_mem_0__127__N_6752[11]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [11])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i12.GSR = "ENABLED";
    FD1P3AX key_mem_14___i13 (.D(key_mem_0__127__N_6752[12]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [12])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i13.GSR = "ENABLED";
    FD1P3AX key_mem_14___i14 (.D(key_mem_0__127__N_6752[13]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [13])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i14.GSR = "ENABLED";
    FD1P3AX key_mem_14___i15 (.D(key_mem_0__127__N_6752[14]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [14])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i15.GSR = "ENABLED";
    FD1P3AX key_mem_14___i16 (.D(key_mem_0__127__N_6752[15]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [15])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i16.GSR = "ENABLED";
    FD1P3AX key_mem_14___i17 (.D(key_mem_0__127__N_6752[16]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [16])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i17.GSR = "ENABLED";
    FD1P3AX key_mem_14___i18 (.D(key_mem_0__127__N_6752[17]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [17])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i18.GSR = "ENABLED";
    FD1P3AX key_mem_14___i19 (.D(key_mem_0__127__N_6752[18]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [18])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i19.GSR = "ENABLED";
    FD1P3AX key_mem_14___i20 (.D(key_mem_0__127__N_6752[19]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [19])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i20.GSR = "ENABLED";
    FD1P3AX key_mem_14___i21 (.D(key_mem_0__127__N_6752[20]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [20])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i21.GSR = "ENABLED";
    FD1P3AX key_mem_14___i22 (.D(key_mem_0__127__N_6752[21]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [21])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i22.GSR = "ENABLED";
    FD1P3AX key_mem_14___i23 (.D(key_mem_0__127__N_6752[22]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [22])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i23.GSR = "ENABLED";
    FD1P3AX key_mem_14___i24 (.D(key_mem_0__127__N_6752[23]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [23])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i24.GSR = "ENABLED";
    FD1P3AX key_mem_14___i25 (.D(key_mem_0__127__N_6752[24]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [24])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i25.GSR = "ENABLED";
    FD1P3AX key_mem_14___i26 (.D(key_mem_0__127__N_6752[25]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [25])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i26.GSR = "ENABLED";
    FD1P3AX key_mem_14___i27 (.D(key_mem_0__127__N_6752[26]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [26])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i27.GSR = "ENABLED";
    FD1P3AX key_mem_14___i28 (.D(key_mem_0__127__N_6752[27]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [27])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i28.GSR = "ENABLED";
    FD1P3AX key_mem_14___i29 (.D(key_mem_0__127__N_6752[28]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [28])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i29.GSR = "ENABLED";
    FD1P3AX key_mem_14___i30 (.D(key_mem_0__127__N_6752[29]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [29])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i30.GSR = "ENABLED";
    FD1P3AX key_mem_14___i31 (.D(key_mem_0__127__N_6752[30]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [30])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i31.GSR = "ENABLED";
    FD1P3AX key_mem_14___i32 (.D(key_mem_0__127__N_6752[31]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [31])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i32.GSR = "ENABLED";
    FD1P3AX key_mem_14___i33 (.D(key_mem_0__127__N_6752[32]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [32])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i33.GSR = "ENABLED";
    FD1P3AX key_mem_14___i34 (.D(key_mem_0__127__N_6752[33]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [33])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i34.GSR = "ENABLED";
    FD1P3AX key_mem_14___i35 (.D(key_mem_0__127__N_6752[34]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [34])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i35.GSR = "ENABLED";
    FD1P3AX key_mem_14___i36 (.D(key_mem_0__127__N_6752[35]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [35])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i36.GSR = "ENABLED";
    FD1P3AX key_mem_14___i37 (.D(key_mem_0__127__N_6752[36]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [36])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i37.GSR = "ENABLED";
    FD1P3AX key_mem_14___i38 (.D(key_mem_0__127__N_6752[37]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [37])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i38.GSR = "ENABLED";
    FD1P3AX key_mem_14___i39 (.D(key_mem_0__127__N_6752[38]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [38])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i39.GSR = "ENABLED";
    FD1P3AX key_mem_14___i40 (.D(key_mem_0__127__N_6752[39]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [39])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i40.GSR = "ENABLED";
    FD1P3AX key_mem_14___i41 (.D(key_mem_0__127__N_6752[40]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [40])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i41.GSR = "ENABLED";
    FD1P3AX key_mem_14___i42 (.D(key_mem_0__127__N_6752[41]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [41])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i42.GSR = "ENABLED";
    FD1P3AX key_mem_14___i43 (.D(key_mem_0__127__N_6752[42]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [42])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i43.GSR = "ENABLED";
    FD1P3AX key_mem_14___i44 (.D(key_mem_0__127__N_6752[43]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [43])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i44.GSR = "ENABLED";
    FD1P3AX key_mem_14___i45 (.D(key_mem_0__127__N_6752[44]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [44])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i45.GSR = "ENABLED";
    FD1P3AX key_mem_14___i46 (.D(key_mem_0__127__N_6752[45]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [45])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i46.GSR = "ENABLED";
    FD1P3AX key_mem_14___i47 (.D(key_mem_0__127__N_6752[46]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [46])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i47.GSR = "ENABLED";
    FD1P3AX key_mem_14___i48 (.D(key_mem_0__127__N_6752[47]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [47])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i48.GSR = "ENABLED";
    FD1P3AX key_mem_14___i49 (.D(key_mem_0__127__N_6752[48]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [48])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i49.GSR = "ENABLED";
    FD1P3AX key_mem_14___i50 (.D(key_mem_0__127__N_6752[49]), .SP(clk_c_enable_436), 
            .CK(clk_c), .Q(\key_mem[14] [49])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i50.GSR = "ENABLED";
    FD1P3AX key_mem_14___i51 (.D(key_mem_0__127__N_6752[50]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [50])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i51.GSR = "ENABLED";
    FD1P3AX key_mem_14___i52 (.D(key_mem_0__127__N_6752[51]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [51])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i52.GSR = "ENABLED";
    FD1P3AX key_mem_14___i53 (.D(key_mem_0__127__N_6752[52]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [52])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i53.GSR = "ENABLED";
    FD1P3AX key_mem_14___i54 (.D(key_mem_0__127__N_6752[53]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [53])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i54.GSR = "ENABLED";
    FD1P3AX key_mem_14___i55 (.D(key_mem_0__127__N_6752[54]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [54])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i55.GSR = "ENABLED";
    FD1P3AX key_mem_14___i56 (.D(key_mem_0__127__N_6752[55]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [55])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i56.GSR = "ENABLED";
    FD1P3AX key_mem_14___i57 (.D(key_mem_0__127__N_6752[56]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [56])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i57.GSR = "ENABLED";
    FD1P3AX key_mem_14___i58 (.D(key_mem_0__127__N_6752[57]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [57])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i58.GSR = "ENABLED";
    FD1P3AX key_mem_14___i59 (.D(key_mem_0__127__N_6752[58]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [58])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i59.GSR = "ENABLED";
    FD1P3AX key_mem_14___i60 (.D(key_mem_0__127__N_6752[59]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [59])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i60.GSR = "ENABLED";
    FD1P3AX key_mem_14___i61 (.D(key_mem_0__127__N_6752[60]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [60])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i61.GSR = "ENABLED";
    FD1P3AX key_mem_14___i62 (.D(key_mem_0__127__N_6752[61]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [61])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i62.GSR = "ENABLED";
    FD1P3AX key_mem_14___i63 (.D(key_mem_0__127__N_6752[62]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [62])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i63.GSR = "ENABLED";
    FD1P3AX key_mem_14___i64 (.D(key_mem_0__127__N_6752[63]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [63])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i64.GSR = "ENABLED";
    FD1P3AX key_mem_14___i65 (.D(key_mem_0__127__N_6752[64]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [64])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i65.GSR = "ENABLED";
    FD1P3AX key_mem_14___i66 (.D(key_mem_0__127__N_6752[65]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [65])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i66.GSR = "ENABLED";
    FD1P3AX key_mem_14___i67 (.D(key_mem_0__127__N_6752[66]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [66])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i67.GSR = "ENABLED";
    FD1P3AX key_mem_14___i68 (.D(key_mem_0__127__N_6752[67]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [67])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i68.GSR = "ENABLED";
    FD1P3AX key_mem_14___i69 (.D(key_mem_0__127__N_6752[68]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [68])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i69.GSR = "ENABLED";
    FD1P3AX key_mem_14___i70 (.D(key_mem_0__127__N_6752[69]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [69])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i70.GSR = "ENABLED";
    FD1P3AX key_mem_14___i71 (.D(key_mem_0__127__N_6752[70]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [70])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i71.GSR = "ENABLED";
    FD1P3AX key_mem_14___i72 (.D(key_mem_0__127__N_6752[71]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [71])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i72.GSR = "ENABLED";
    FD1P3AX key_mem_14___i73 (.D(key_mem_0__127__N_6752[72]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [72])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i73.GSR = "ENABLED";
    FD1P3AX key_mem_14___i74 (.D(key_mem_0__127__N_6752[73]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [73])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i74.GSR = "ENABLED";
    FD1P3AX key_mem_14___i75 (.D(key_mem_0__127__N_6752[74]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [74])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i75.GSR = "ENABLED";
    FD1P3AX key_mem_14___i76 (.D(key_mem_0__127__N_6752[75]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [75])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i76.GSR = "ENABLED";
    FD1P3AX key_mem_14___i77 (.D(key_mem_0__127__N_6752[76]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [76])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i77.GSR = "ENABLED";
    FD1P3AX key_mem_14___i78 (.D(key_mem_0__127__N_6752[77]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [77])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i78.GSR = "ENABLED";
    FD1P3AX key_mem_14___i79 (.D(key_mem_0__127__N_6752[78]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [78])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i79.GSR = "ENABLED";
    FD1P3AX key_mem_14___i80 (.D(key_mem_0__127__N_6752[79]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [79])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i80.GSR = "ENABLED";
    FD1P3AX key_mem_14___i81 (.D(key_mem_0__127__N_6752[80]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [80])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i81.GSR = "ENABLED";
    FD1P3AX key_mem_14___i82 (.D(key_mem_0__127__N_6752[81]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [81])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i82.GSR = "ENABLED";
    FD1P3AX key_mem_14___i83 (.D(key_mem_0__127__N_6752[82]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [82])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i83.GSR = "ENABLED";
    FD1P3AX key_mem_14___i84 (.D(key_mem_0__127__N_6752[83]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [83])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i84.GSR = "ENABLED";
    FD1P3AX key_mem_14___i85 (.D(key_mem_0__127__N_6752[84]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [84])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i85.GSR = "ENABLED";
    FD1P3AX key_mem_14___i86 (.D(key_mem_0__127__N_6752[85]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [85])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i86.GSR = "ENABLED";
    FD1P3AX key_mem_14___i87 (.D(key_mem_0__127__N_6752[86]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [86])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i87.GSR = "ENABLED";
    FD1P3AX key_mem_14___i88 (.D(key_mem_0__127__N_6752[87]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [87])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i88.GSR = "ENABLED";
    FD1P3AX key_mem_14___i89 (.D(key_mem_0__127__N_6752[88]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [88])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i89.GSR = "ENABLED";
    FD1P3AX key_mem_14___i90 (.D(key_mem_0__127__N_6752[89]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [89])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i90.GSR = "ENABLED";
    FD1P3AX key_mem_14___i91 (.D(key_mem_0__127__N_6752[90]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [90])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i91.GSR = "ENABLED";
    FD1P3AX key_mem_14___i92 (.D(key_mem_0__127__N_6752[91]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [91])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i92.GSR = "ENABLED";
    FD1P3AX key_mem_14___i93 (.D(key_mem_0__127__N_6752[92]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [92])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i93.GSR = "ENABLED";
    FD1P3AX key_mem_14___i94 (.D(key_mem_0__127__N_6752[93]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [93])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i94.GSR = "ENABLED";
    FD1P3AX key_mem_14___i95 (.D(key_mem_0__127__N_6752[94]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [94])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i95.GSR = "ENABLED";
    FD1P3AX key_mem_14___i96 (.D(key_mem_0__127__N_6752[95]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [95])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i96.GSR = "ENABLED";
    FD1P3AX key_mem_14___i97 (.D(key_mem_0__127__N_6752[96]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [96])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i97.GSR = "ENABLED";
    FD1P3AX key_mem_14___i98 (.D(key_mem_0__127__N_6752[97]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [97])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i98.GSR = "ENABLED";
    FD1P3AX key_mem_14___i99 (.D(key_mem_0__127__N_6752[98]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [98])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i99.GSR = "ENABLED";
    FD1P3AX key_mem_14___i100 (.D(key_mem_0__127__N_6752[99]), .SP(clk_c_enable_486), 
            .CK(clk_c), .Q(\key_mem[14] [99])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i100.GSR = "ENABLED";
    FD1P3AX key_mem_14___i101 (.D(key_mem_0__127__N_6752[100]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[14] [100])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i101.GSR = "ENABLED";
    FD1P3AX key_mem_14___i102 (.D(key_mem_0__127__N_6752[101]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[14] [101])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i102.GSR = "ENABLED";
    FD1P3AX key_mem_14___i103 (.D(key_mem_0__127__N_6752[102]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[14] [102])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i103.GSR = "ENABLED";
    FD1P3AX key_mem_14___i104 (.D(key_mem_0__127__N_6752[103]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[14] [103])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i104.GSR = "ENABLED";
    FD1P3AX key_mem_14___i105 (.D(key_mem_0__127__N_6752[104]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[14] [104])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i105.GSR = "ENABLED";
    FD1P3AX key_mem_14___i106 (.D(key_mem_0__127__N_6752[105]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[14] [105])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i106.GSR = "ENABLED";
    FD1P3AX key_mem_14___i107 (.D(key_mem_0__127__N_6752[106]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[14] [106])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i107.GSR = "ENABLED";
    FD1P3AX key_mem_14___i108 (.D(key_mem_0__127__N_6752[107]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[14] [107])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i108.GSR = "ENABLED";
    FD1P3AX key_mem_14___i109 (.D(key_mem_0__127__N_6752[108]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[14] [108])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i109.GSR = "ENABLED";
    FD1P3AX key_mem_14___i110 (.D(key_mem_0__127__N_6752[109]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[14] [109])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i110.GSR = "ENABLED";
    FD1P3AX key_mem_14___i111 (.D(key_mem_0__127__N_6752[110]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[14] [110])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i111.GSR = "ENABLED";
    FD1P3AX key_mem_14___i112 (.D(key_mem_0__127__N_6752[111]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[14] [111])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i112.GSR = "ENABLED";
    FD1P3AX key_mem_14___i113 (.D(key_mem_0__127__N_6752[112]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[14] [112])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i113.GSR = "ENABLED";
    FD1P3AX key_mem_14___i114 (.D(key_mem_0__127__N_6752[113]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[14] [113])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i114.GSR = "ENABLED";
    FD1P3AX key_mem_14___i115 (.D(key_mem_0__127__N_6752[114]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[14] [114])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i115.GSR = "ENABLED";
    FD1P3AX key_mem_14___i116 (.D(key_mem_0__127__N_6752[115]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[14] [115])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i116.GSR = "ENABLED";
    FD1P3AX key_mem_14___i117 (.D(key_mem_0__127__N_6752[116]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[14] [116])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i117.GSR = "ENABLED";
    FD1P3AX key_mem_14___i118 (.D(key_mem_0__127__N_6752[117]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[14] [117])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i118.GSR = "ENABLED";
    FD1P3AX key_mem_14___i119 (.D(key_mem_0__127__N_6752[118]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[14] [118])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i119.GSR = "ENABLED";
    FD1P3AX key_mem_14___i120 (.D(key_mem_0__127__N_6752[119]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[14] [119])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i120.GSR = "ENABLED";
    FD1P3AX key_mem_14___i121 (.D(key_mem_0__127__N_6752[120]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[14] [120])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i121.GSR = "ENABLED";
    FD1P3AX key_mem_14___i122 (.D(key_mem_0__127__N_6752[121]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[14] [121])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i122.GSR = "ENABLED";
    FD1P3AX key_mem_14___i123 (.D(key_mem_0__127__N_6752[122]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[14] [122])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i123.GSR = "ENABLED";
    FD1P3AX key_mem_14___i124 (.D(key_mem_0__127__N_6752[123]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[14] [123])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i124.GSR = "ENABLED";
    FD1P3AX key_mem_14___i125 (.D(key_mem_0__127__N_6752[124]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[14] [124])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i125.GSR = "ENABLED";
    FD1P3AX key_mem_14___i126 (.D(key_mem_0__127__N_6752[125]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[14] [125])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i126.GSR = "ENABLED";
    FD1P3AX key_mem_14___i127 (.D(key_mem_0__127__N_6752[126]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[14] [126])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i127.GSR = "ENABLED";
    FD1P3AX key_mem_14___i128 (.D(key_mem_0__127__N_6752[127]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[14] [127])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i128.GSR = "ENABLED";
    FD1P3AX key_mem_14___i129 (.D(key_mem_0__127__N_6624[0]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[13] [0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i129.GSR = "ENABLED";
    FD1P3AX key_mem_14___i130 (.D(key_mem_0__127__N_6624[1]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[13] [1])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i130.GSR = "ENABLED";
    FD1P3AX key_mem_14___i131 (.D(key_mem_0__127__N_6624[2]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[13] [2])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i131.GSR = "ENABLED";
    FD1P3AX key_mem_14___i132 (.D(key_mem_0__127__N_6624[3]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[13] [3])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i132.GSR = "ENABLED";
    FD1P3AX key_mem_14___i133 (.D(key_mem_0__127__N_6624[4]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[13] [4])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i133.GSR = "ENABLED";
    FD1P3AX key_mem_14___i134 (.D(key_mem_0__127__N_6624[5]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[13] [5])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i134.GSR = "ENABLED";
    FD1P3AX key_mem_14___i135 (.D(key_mem_0__127__N_6624[6]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[13] [6])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i135.GSR = "ENABLED";
    FD1P3AX key_mem_14___i136 (.D(key_mem_0__127__N_6624[7]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[13] [7])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i136.GSR = "ENABLED";
    FD1P3AX key_mem_14___i137 (.D(key_mem_0__127__N_6624[8]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[13] [8])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i137.GSR = "ENABLED";
    FD1P3AX key_mem_14___i138 (.D(key_mem_0__127__N_6624[9]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[13] [9])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i138.GSR = "ENABLED";
    FD1P3AX key_mem_14___i139 (.D(key_mem_0__127__N_6624[10]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[13] [10])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i139.GSR = "ENABLED";
    FD1P3AX key_mem_14___i140 (.D(key_mem_0__127__N_6624[11]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[13] [11])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i140.GSR = "ENABLED";
    FD1P3AX key_mem_14___i141 (.D(key_mem_0__127__N_6624[12]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[13] [12])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i141.GSR = "ENABLED";
    FD1P3AX key_mem_14___i142 (.D(key_mem_0__127__N_6624[13]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[13] [13])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i142.GSR = "ENABLED";
    FD1P3AX key_mem_14___i143 (.D(key_mem_0__127__N_6624[14]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[13] [14])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i143.GSR = "ENABLED";
    FD1P3AX key_mem_14___i144 (.D(key_mem_0__127__N_6624[15]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[13] [15])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i144.GSR = "ENABLED";
    FD1P3AX key_mem_14___i145 (.D(key_mem_0__127__N_6624[16]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[13] [16])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i145.GSR = "ENABLED";
    FD1P3AX key_mem_14___i146 (.D(key_mem_0__127__N_6624[17]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[13] [17])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i146.GSR = "ENABLED";
    FD1P3AX key_mem_14___i147 (.D(key_mem_0__127__N_6624[18]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[13] [18])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i147.GSR = "ENABLED";
    FD1P3AX key_mem_14___i148 (.D(key_mem_0__127__N_6624[19]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[13] [19])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i148.GSR = "ENABLED";
    FD1P3AX key_mem_14___i149 (.D(key_mem_0__127__N_6624[20]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[13] [20])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i149.GSR = "ENABLED";
    FD1P3AX key_mem_14___i150 (.D(key_mem_0__127__N_6624[21]), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(\key_mem[13] [21])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i150.GSR = "ENABLED";
    FD1P3AX key_mem_14___i151 (.D(key_mem_0__127__N_6624[22]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [22])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i151.GSR = "ENABLED";
    FD1P3AX key_mem_14___i152 (.D(key_mem_0__127__N_6624[23]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [23])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i152.GSR = "ENABLED";
    FD1P3AX key_mem_14___i153 (.D(key_mem_0__127__N_6624[24]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [24])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i153.GSR = "ENABLED";
    FD1P3AX key_mem_14___i154 (.D(key_mem_0__127__N_6624[25]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [25])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i154.GSR = "ENABLED";
    FD1P3AX key_mem_14___i155 (.D(key_mem_0__127__N_6624[26]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [26])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i155.GSR = "ENABLED";
    FD1P3AX key_mem_14___i156 (.D(key_mem_0__127__N_6624[27]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [27])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i156.GSR = "ENABLED";
    FD1P3AX key_mem_14___i157 (.D(key_mem_0__127__N_6624[28]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [28])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i157.GSR = "ENABLED";
    FD1P3AX key_mem_14___i158 (.D(key_mem_0__127__N_6624[29]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [29])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i158.GSR = "ENABLED";
    FD1P3AX key_mem_14___i159 (.D(key_mem_0__127__N_6624[30]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [30])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i159.GSR = "ENABLED";
    FD1P3AX key_mem_14___i160 (.D(key_mem_0__127__N_6624[31]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [31])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i160.GSR = "ENABLED";
    FD1P3AX key_mem_14___i161 (.D(key_mem_0__127__N_6624[32]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [32])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i161.GSR = "ENABLED";
    FD1P3AX key_mem_14___i162 (.D(key_mem_0__127__N_6624[33]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [33])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i162.GSR = "ENABLED";
    FD1P3AX key_mem_14___i163 (.D(key_mem_0__127__N_6624[34]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [34])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i163.GSR = "ENABLED";
    FD1P3AX key_mem_14___i164 (.D(key_mem_0__127__N_6624[35]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [35])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i164.GSR = "ENABLED";
    FD1P3AX key_mem_14___i165 (.D(key_mem_0__127__N_6624[36]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [36])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i165.GSR = "ENABLED";
    FD1P3AX key_mem_14___i166 (.D(key_mem_0__127__N_6624[37]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [37])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i166.GSR = "ENABLED";
    FD1P3AX key_mem_14___i167 (.D(key_mem_0__127__N_6624[38]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [38])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i167.GSR = "ENABLED";
    FD1P3AX key_mem_14___i168 (.D(key_mem_0__127__N_6624[39]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [39])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i168.GSR = "ENABLED";
    FD1P3AX key_mem_14___i169 (.D(key_mem_0__127__N_6624[40]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [40])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i169.GSR = "ENABLED";
    FD1P3AX key_mem_14___i170 (.D(key_mem_0__127__N_6624[41]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [41])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i170.GSR = "ENABLED";
    FD1P3AX key_mem_14___i171 (.D(key_mem_0__127__N_6624[42]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [42])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i171.GSR = "ENABLED";
    FD1P3AX key_mem_14___i172 (.D(key_mem_0__127__N_6624[43]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [43])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i172.GSR = "ENABLED";
    FD1P3AX key_mem_14___i173 (.D(key_mem_0__127__N_6624[44]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [44])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i173.GSR = "ENABLED";
    FD1P3AX key_mem_14___i174 (.D(key_mem_0__127__N_6624[45]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [45])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i174.GSR = "ENABLED";
    FD1P3AX key_mem_14___i175 (.D(key_mem_0__127__N_6624[46]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [46])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i175.GSR = "ENABLED";
    FD1P3AX key_mem_14___i176 (.D(key_mem_0__127__N_6624[47]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [47])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i176.GSR = "ENABLED";
    FD1P3AX key_mem_14___i177 (.D(key_mem_0__127__N_6624[48]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [48])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i177.GSR = "ENABLED";
    FD1P3AX key_mem_14___i178 (.D(key_mem_0__127__N_6624[49]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [49])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i178.GSR = "ENABLED";
    FD1P3AX key_mem_14___i179 (.D(key_mem_0__127__N_6624[50]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [50])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i179.GSR = "ENABLED";
    FD1P3AX key_mem_14___i180 (.D(key_mem_0__127__N_6624[51]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [51])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i180.GSR = "ENABLED";
    FD1P3AX key_mem_14___i181 (.D(key_mem_0__127__N_6624[52]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [52])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i181.GSR = "ENABLED";
    FD1P3AX key_mem_14___i182 (.D(key_mem_0__127__N_6624[53]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [53])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i182.GSR = "ENABLED";
    FD1P3AX key_mem_14___i183 (.D(key_mem_0__127__N_6624[54]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [54])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i183.GSR = "ENABLED";
    FD1P3AX key_mem_14___i184 (.D(key_mem_0__127__N_6624[55]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [55])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i184.GSR = "ENABLED";
    FD1P3AX key_mem_14___i185 (.D(key_mem_0__127__N_6624[56]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [56])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i185.GSR = "ENABLED";
    FD1P3AX key_mem_14___i186 (.D(key_mem_0__127__N_6624[57]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [57])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i186.GSR = "ENABLED";
    FD1P3AX key_mem_14___i187 (.D(key_mem_0__127__N_6624[58]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [58])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i187.GSR = "ENABLED";
    FD1P3AX key_mem_14___i188 (.D(key_mem_0__127__N_6624[59]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [59])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i188.GSR = "ENABLED";
    FD1P3AX key_mem_14___i189 (.D(key_mem_0__127__N_6624[60]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [60])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i189.GSR = "ENABLED";
    FD1P3AX key_mem_14___i190 (.D(key_mem_0__127__N_6624[61]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [61])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i190.GSR = "ENABLED";
    FD1P3AX key_mem_14___i191 (.D(key_mem_0__127__N_6624[62]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [62])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i191.GSR = "ENABLED";
    FD1P3AX key_mem_14___i192 (.D(key_mem_0__127__N_6624[63]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [63])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i192.GSR = "ENABLED";
    FD1P3AX key_mem_14___i193 (.D(key_mem_0__127__N_6624[64]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [64])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i193.GSR = "ENABLED";
    FD1P3AX key_mem_14___i194 (.D(key_mem_0__127__N_6624[65]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [65])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i194.GSR = "ENABLED";
    FD1P3AX key_mem_14___i195 (.D(key_mem_0__127__N_6624[66]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [66])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i195.GSR = "ENABLED";
    FD1P3AX key_mem_14___i196 (.D(key_mem_0__127__N_6624[67]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [67])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i196.GSR = "ENABLED";
    FD1P3AX key_mem_14___i197 (.D(key_mem_0__127__N_6624[68]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [68])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i197.GSR = "ENABLED";
    FD1P3AX key_mem_14___i198 (.D(key_mem_0__127__N_6624[69]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [69])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i198.GSR = "ENABLED";
    FD1P3AX key_mem_14___i199 (.D(key_mem_0__127__N_6624[70]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [70])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i199.GSR = "ENABLED";
    FD1P3AX key_mem_14___i200 (.D(key_mem_0__127__N_6624[71]), .SP(clk_c_enable_586), 
            .CK(clk_c), .Q(\key_mem[13] [71])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i200.GSR = "ENABLED";
    FD1P3AX key_mem_14___i201 (.D(key_mem_0__127__N_6624[72]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [72])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i201.GSR = "ENABLED";
    FD1P3AX key_mem_14___i202 (.D(key_mem_0__127__N_6624[73]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [73])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i202.GSR = "ENABLED";
    FD1P3AX key_mem_14___i203 (.D(key_mem_0__127__N_6624[74]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [74])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i203.GSR = "ENABLED";
    FD1P3AX key_mem_14___i204 (.D(key_mem_0__127__N_6624[75]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [75])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i204.GSR = "ENABLED";
    FD1P3AX key_mem_14___i205 (.D(key_mem_0__127__N_6624[76]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [76])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i205.GSR = "ENABLED";
    FD1P3AX key_mem_14___i206 (.D(key_mem_0__127__N_6624[77]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [77])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i206.GSR = "ENABLED";
    FD1P3AX key_mem_14___i207 (.D(key_mem_0__127__N_6624[78]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [78])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i207.GSR = "ENABLED";
    FD1P3AX key_mem_14___i208 (.D(key_mem_0__127__N_6624[79]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [79])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i208.GSR = "ENABLED";
    FD1P3AX key_mem_14___i209 (.D(key_mem_0__127__N_6624[80]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [80])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i209.GSR = "ENABLED";
    FD1P3AX key_mem_14___i210 (.D(key_mem_0__127__N_6624[81]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [81])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i210.GSR = "ENABLED";
    FD1P3AX key_mem_14___i211 (.D(key_mem_0__127__N_6624[82]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [82])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i211.GSR = "ENABLED";
    FD1P3AX key_mem_14___i212 (.D(key_mem_0__127__N_6624[83]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [83])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i212.GSR = "ENABLED";
    FD1P3AX key_mem_14___i213 (.D(key_mem_0__127__N_6624[84]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [84])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i213.GSR = "ENABLED";
    FD1P3AX key_mem_14___i214 (.D(key_mem_0__127__N_6624[85]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [85])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i214.GSR = "ENABLED";
    FD1P3AX key_mem_14___i215 (.D(key_mem_0__127__N_6624[86]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [86])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i215.GSR = "ENABLED";
    FD1P3AX key_mem_14___i216 (.D(key_mem_0__127__N_6624[87]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [87])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i216.GSR = "ENABLED";
    FD1P3AX key_mem_14___i217 (.D(key_mem_0__127__N_6624[88]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [88])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i217.GSR = "ENABLED";
    FD1P3AX key_mem_14___i218 (.D(key_mem_0__127__N_6624[89]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [89])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i218.GSR = "ENABLED";
    FD1P3AX key_mem_14___i219 (.D(key_mem_0__127__N_6624[90]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [90])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i219.GSR = "ENABLED";
    FD1P3AX key_mem_14___i220 (.D(key_mem_0__127__N_6624[91]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [91])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i220.GSR = "ENABLED";
    FD1P3AX key_mem_14___i221 (.D(key_mem_0__127__N_6624[92]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [92])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i221.GSR = "ENABLED";
    FD1P3AX key_mem_14___i222 (.D(key_mem_0__127__N_6624[93]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [93])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i222.GSR = "ENABLED";
    FD1P3AX key_mem_14___i223 (.D(key_mem_0__127__N_6624[94]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [94])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i223.GSR = "ENABLED";
    FD1P3AX key_mem_14___i224 (.D(key_mem_0__127__N_6624[95]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [95])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i224.GSR = "ENABLED";
    FD1P3AX key_mem_14___i225 (.D(key_mem_0__127__N_6624[96]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [96])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i225.GSR = "ENABLED";
    FD1P3AX key_mem_14___i226 (.D(key_mem_0__127__N_6624[97]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [97])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i226.GSR = "ENABLED";
    FD1P3AX key_mem_14___i227 (.D(key_mem_0__127__N_6624[98]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [98])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i227.GSR = "ENABLED";
    FD1P3AX key_mem_14___i228 (.D(key_mem_0__127__N_6624[99]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [99])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i228.GSR = "ENABLED";
    FD1P3AX key_mem_14___i229 (.D(key_mem_0__127__N_6624[100]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [100])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i229.GSR = "ENABLED";
    FD1P3AX key_mem_14___i230 (.D(key_mem_0__127__N_6624[101]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [101])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i230.GSR = "ENABLED";
    FD1P3AX key_mem_14___i231 (.D(key_mem_0__127__N_6624[102]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [102])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i231.GSR = "ENABLED";
    FD1P3AX key_mem_14___i232 (.D(key_mem_0__127__N_6624[103]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [103])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i232.GSR = "ENABLED";
    FD1P3AX key_mem_14___i233 (.D(key_mem_0__127__N_6624[104]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [104])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i233.GSR = "ENABLED";
    FD1P3AX key_mem_14___i234 (.D(key_mem_0__127__N_6624[105]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [105])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i234.GSR = "ENABLED";
    FD1P3AX key_mem_14___i235 (.D(key_mem_0__127__N_6624[106]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [106])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i235.GSR = "ENABLED";
    FD1P3AX key_mem_14___i236 (.D(key_mem_0__127__N_6624[107]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [107])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i236.GSR = "ENABLED";
    FD1P3AX key_mem_14___i237 (.D(key_mem_0__127__N_6624[108]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [108])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i237.GSR = "ENABLED";
    FD1P3AX key_mem_14___i238 (.D(key_mem_0__127__N_6624[109]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [109])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i238.GSR = "ENABLED";
    FD1P3AX key_mem_14___i239 (.D(key_mem_0__127__N_6624[110]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [110])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i239.GSR = "ENABLED";
    FD1P3AX key_mem_14___i240 (.D(key_mem_0__127__N_6624[111]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [111])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i240.GSR = "ENABLED";
    FD1P3AX key_mem_14___i241 (.D(key_mem_0__127__N_6624[112]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [112])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i241.GSR = "ENABLED";
    FD1P3AX key_mem_14___i242 (.D(key_mem_0__127__N_6624[113]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [113])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i242.GSR = "ENABLED";
    FD1P3AX key_mem_14___i243 (.D(key_mem_0__127__N_6624[114]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [114])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i243.GSR = "ENABLED";
    FD1P3AX key_mem_14___i244 (.D(key_mem_0__127__N_6624[115]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [115])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i244.GSR = "ENABLED";
    FD1P3AX key_mem_14___i245 (.D(key_mem_0__127__N_6624[116]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [116])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i245.GSR = "ENABLED";
    FD1P3AX key_mem_14___i246 (.D(key_mem_0__127__N_6624[117]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [117])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i246.GSR = "ENABLED";
    FD1P3AX key_mem_14___i247 (.D(key_mem_0__127__N_6624[118]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [118])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i247.GSR = "ENABLED";
    FD1P3AX key_mem_14___i248 (.D(key_mem_0__127__N_6624[119]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [119])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i248.GSR = "ENABLED";
    FD1P3AX key_mem_14___i249 (.D(key_mem_0__127__N_6624[120]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [120])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i249.GSR = "ENABLED";
    FD1P3AX key_mem_14___i250 (.D(key_mem_0__127__N_6624[121]), .SP(clk_c_enable_636), 
            .CK(clk_c), .Q(\key_mem[13] [121])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i250.GSR = "ENABLED";
    FD1P3AX key_mem_14___i251 (.D(key_mem_0__127__N_6624[122]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[13] [122])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i251.GSR = "ENABLED";
    FD1P3AX key_mem_14___i252 (.D(key_mem_0__127__N_6624[123]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[13] [123])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i252.GSR = "ENABLED";
    FD1P3AX key_mem_14___i253 (.D(key_mem_0__127__N_6624[124]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[13] [124])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i253.GSR = "ENABLED";
    FD1P3AX key_mem_14___i254 (.D(key_mem_0__127__N_6624[125]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[13] [125])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i254.GSR = "ENABLED";
    FD1P3AX key_mem_14___i255 (.D(key_mem_0__127__N_6624[126]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[13] [126])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i255.GSR = "ENABLED";
    FD1P3AX key_mem_14___i256 (.D(key_mem_0__127__N_6624[127]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[13] [127])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i256.GSR = "ENABLED";
    FD1P3AX key_mem_14___i257 (.D(key_mem_0__127__N_6496[0]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[12] [0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i257.GSR = "ENABLED";
    FD1P3AX key_mem_14___i258 (.D(key_mem_0__127__N_6496[1]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[12] [1])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i258.GSR = "ENABLED";
    FD1P3AX key_mem_14___i259 (.D(key_mem_0__127__N_6496[2]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[12] [2])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i259.GSR = "ENABLED";
    FD1P3AX key_mem_14___i260 (.D(key_mem_0__127__N_6496[3]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[12] [3])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i260.GSR = "ENABLED";
    FD1P3AX key_mem_14___i261 (.D(key_mem_0__127__N_6496[4]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[12] [4])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i261.GSR = "ENABLED";
    FD1P3AX key_mem_14___i262 (.D(key_mem_0__127__N_6496[5]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[12] [5])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i262.GSR = "ENABLED";
    FD1P3AX key_mem_14___i263 (.D(key_mem_0__127__N_6496[6]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[12] [6])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i263.GSR = "ENABLED";
    FD1P3AX key_mem_14___i264 (.D(key_mem_0__127__N_6496[7]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[12] [7])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i264.GSR = "ENABLED";
    FD1P3AX key_mem_14___i265 (.D(key_mem_0__127__N_6496[8]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[12] [8])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i265.GSR = "ENABLED";
    FD1P3AX key_mem_14___i266 (.D(key_mem_0__127__N_6496[9]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[12] [9])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i266.GSR = "ENABLED";
    FD1P3AX key_mem_14___i267 (.D(key_mem_0__127__N_6496[10]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[12] [10])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i267.GSR = "ENABLED";
    FD1P3AX key_mem_14___i268 (.D(key_mem_0__127__N_6496[11]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[12] [11])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i268.GSR = "ENABLED";
    FD1P3AX key_mem_14___i269 (.D(key_mem_0__127__N_6496[12]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[12] [12])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i269.GSR = "ENABLED";
    FD1P3AX key_mem_14___i270 (.D(key_mem_0__127__N_6496[13]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[12] [13])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i270.GSR = "ENABLED";
    FD1P3AX key_mem_14___i271 (.D(key_mem_0__127__N_6496[14]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[12] [14])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i271.GSR = "ENABLED";
    FD1P3AX key_mem_14___i272 (.D(key_mem_0__127__N_6496[15]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[12] [15])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i272.GSR = "ENABLED";
    FD1P3AX key_mem_14___i273 (.D(key_mem_0__127__N_6496[16]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[12] [16])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i273.GSR = "ENABLED";
    FD1P3AX key_mem_14___i274 (.D(key_mem_0__127__N_6496[17]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[12] [17])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i274.GSR = "ENABLED";
    FD1P3AX key_mem_14___i275 (.D(key_mem_0__127__N_6496[18]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[12] [18])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i275.GSR = "ENABLED";
    FD1P3AX key_mem_14___i276 (.D(key_mem_0__127__N_6496[19]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[12] [19])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i276.GSR = "ENABLED";
    FD1P3AX key_mem_14___i277 (.D(key_mem_0__127__N_6496[20]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[12] [20])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i277.GSR = "ENABLED";
    FD1P3AX key_mem_14___i278 (.D(key_mem_0__127__N_6496[21]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[12] [21])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i278.GSR = "ENABLED";
    FD1P3AX key_mem_14___i279 (.D(key_mem_0__127__N_6496[22]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[12] [22])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i279.GSR = "ENABLED";
    FD1P3AX key_mem_14___i280 (.D(key_mem_0__127__N_6496[23]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[12] [23])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i280.GSR = "ENABLED";
    FD1P3AX key_mem_14___i281 (.D(key_mem_0__127__N_6496[24]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[12] [24])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i281.GSR = "ENABLED";
    FD1P3AX key_mem_14___i282 (.D(key_mem_0__127__N_6496[25]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[12] [25])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i282.GSR = "ENABLED";
    FD1P3AX key_mem_14___i283 (.D(key_mem_0__127__N_6496[26]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[12] [26])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i283.GSR = "ENABLED";
    FD1P3AX key_mem_14___i284 (.D(key_mem_0__127__N_6496[27]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[12] [27])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i284.GSR = "ENABLED";
    FD1P3AX key_mem_14___i285 (.D(key_mem_0__127__N_6496[28]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[12] [28])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i285.GSR = "ENABLED";
    FD1P3AX key_mem_14___i286 (.D(key_mem_0__127__N_6496[29]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[12] [29])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i286.GSR = "ENABLED";
    FD1P3AX key_mem_14___i287 (.D(key_mem_0__127__N_6496[30]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[12] [30])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i287.GSR = "ENABLED";
    FD1P3AX key_mem_14___i288 (.D(key_mem_0__127__N_6496[31]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[12] [31])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i288.GSR = "ENABLED";
    FD1P3AX key_mem_14___i289 (.D(key_mem_0__127__N_6496[32]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[12] [32])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i289.GSR = "ENABLED";
    FD1P3AX key_mem_14___i290 (.D(key_mem_0__127__N_6496[33]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[12] [33])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i290.GSR = "ENABLED";
    FD1P3AX key_mem_14___i291 (.D(key_mem_0__127__N_6496[34]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[12] [34])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i291.GSR = "ENABLED";
    FD1P3AX key_mem_14___i292 (.D(key_mem_0__127__N_6496[35]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[12] [35])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i292.GSR = "ENABLED";
    FD1P3AX key_mem_14___i293 (.D(key_mem_0__127__N_6496[36]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[12] [36])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i293.GSR = "ENABLED";
    FD1P3AX key_mem_14___i294 (.D(key_mem_0__127__N_6496[37]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[12] [37])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i294.GSR = "ENABLED";
    FD1P3AX key_mem_14___i295 (.D(key_mem_0__127__N_6496[38]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[12] [38])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i295.GSR = "ENABLED";
    FD1P3AX key_mem_14___i296 (.D(key_mem_0__127__N_6496[39]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[12] [39])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i296.GSR = "ENABLED";
    FD1P3AX key_mem_14___i297 (.D(key_mem_0__127__N_6496[40]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[12] [40])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i297.GSR = "ENABLED";
    FD1P3AX key_mem_14___i298 (.D(key_mem_0__127__N_6496[41]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[12] [41])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i298.GSR = "ENABLED";
    FD1P3AX key_mem_14___i299 (.D(key_mem_0__127__N_6496[42]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[12] [42])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i299.GSR = "ENABLED";
    FD1P3AX key_mem_14___i300 (.D(key_mem_0__127__N_6496[43]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(\key_mem[12] [43])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i300.GSR = "ENABLED";
    FD1P3AX key_mem_14___i301 (.D(key_mem_0__127__N_6496[44]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [44])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i301.GSR = "ENABLED";
    FD1P3AX key_mem_14___i302 (.D(key_mem_0__127__N_6496[45]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [45])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i302.GSR = "ENABLED";
    FD1P3AX key_mem_14___i303 (.D(key_mem_0__127__N_6496[46]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [46])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i303.GSR = "ENABLED";
    FD1P3AX key_mem_14___i304 (.D(key_mem_0__127__N_6496[47]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [47])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i304.GSR = "ENABLED";
    FD1P3AX key_mem_14___i305 (.D(key_mem_0__127__N_6496[48]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [48])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i305.GSR = "ENABLED";
    FD1P3AX key_mem_14___i306 (.D(key_mem_0__127__N_6496[49]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [49])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i306.GSR = "ENABLED";
    FD1P3AX key_mem_14___i307 (.D(key_mem_0__127__N_6496[50]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [50])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i307.GSR = "ENABLED";
    FD1P3AX key_mem_14___i308 (.D(key_mem_0__127__N_6496[51]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [51])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i308.GSR = "ENABLED";
    FD1P3AX key_mem_14___i309 (.D(key_mem_0__127__N_6496[52]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [52])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i309.GSR = "ENABLED";
    FD1P3AX key_mem_14___i310 (.D(key_mem_0__127__N_6496[53]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [53])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i310.GSR = "ENABLED";
    FD1P3AX key_mem_14___i311 (.D(key_mem_0__127__N_6496[54]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [54])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i311.GSR = "ENABLED";
    FD1P3AX key_mem_14___i312 (.D(key_mem_0__127__N_6496[55]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [55])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i312.GSR = "ENABLED";
    FD1P3AX key_mem_14___i313 (.D(key_mem_0__127__N_6496[56]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [56])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i313.GSR = "ENABLED";
    FD1P3AX key_mem_14___i314 (.D(key_mem_0__127__N_6496[57]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [57])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i314.GSR = "ENABLED";
    FD1P3AX key_mem_14___i315 (.D(key_mem_0__127__N_6496[58]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [58])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i315.GSR = "ENABLED";
    FD1P3AX key_mem_14___i316 (.D(key_mem_0__127__N_6496[59]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [59])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i316.GSR = "ENABLED";
    FD1P3AX key_mem_14___i317 (.D(key_mem_0__127__N_6496[60]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [60])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i317.GSR = "ENABLED";
    FD1P3AX key_mem_14___i318 (.D(key_mem_0__127__N_6496[61]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [61])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i318.GSR = "ENABLED";
    FD1P3AX key_mem_14___i319 (.D(key_mem_0__127__N_6496[62]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [62])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i319.GSR = "ENABLED";
    FD1P3AX key_mem_14___i320 (.D(key_mem_0__127__N_6496[63]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [63])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i320.GSR = "ENABLED";
    FD1P3AX key_mem_14___i321 (.D(key_mem_0__127__N_6496[64]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [64])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i321.GSR = "ENABLED";
    FD1P3AX key_mem_14___i322 (.D(key_mem_0__127__N_6496[65]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [65])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i322.GSR = "ENABLED";
    FD1P3AX key_mem_14___i323 (.D(key_mem_0__127__N_6496[66]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [66])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i323.GSR = "ENABLED";
    FD1P3AX key_mem_14___i324 (.D(key_mem_0__127__N_6496[67]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [67])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i324.GSR = "ENABLED";
    FD1P3AX key_mem_14___i325 (.D(key_mem_0__127__N_6496[68]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [68])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i325.GSR = "ENABLED";
    FD1P3AX key_mem_14___i326 (.D(key_mem_0__127__N_6496[69]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [69])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i326.GSR = "ENABLED";
    FD1P3AX key_mem_14___i327 (.D(key_mem_0__127__N_6496[70]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [70])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i327.GSR = "ENABLED";
    FD1P3AX key_mem_14___i328 (.D(key_mem_0__127__N_6496[71]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [71])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i328.GSR = "ENABLED";
    FD1P3AX key_mem_14___i329 (.D(key_mem_0__127__N_6496[72]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [72])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i329.GSR = "ENABLED";
    FD1P3AX key_mem_14___i330 (.D(key_mem_0__127__N_6496[73]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [73])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i330.GSR = "ENABLED";
    FD1P3AX key_mem_14___i331 (.D(key_mem_0__127__N_6496[74]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [74])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i331.GSR = "ENABLED";
    FD1P3AX key_mem_14___i332 (.D(key_mem_0__127__N_6496[75]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [75])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i332.GSR = "ENABLED";
    FD1P3AX key_mem_14___i333 (.D(key_mem_0__127__N_6496[76]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [76])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i333.GSR = "ENABLED";
    FD1P3AX key_mem_14___i334 (.D(key_mem_0__127__N_6496[77]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [77])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i334.GSR = "ENABLED";
    FD1P3AX key_mem_14___i335 (.D(key_mem_0__127__N_6496[78]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [78])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i335.GSR = "ENABLED";
    FD1P3AX key_mem_14___i336 (.D(key_mem_0__127__N_6496[79]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [79])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i336.GSR = "ENABLED";
    FD1P3AX key_mem_14___i337 (.D(key_mem_0__127__N_6496[80]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [80])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i337.GSR = "ENABLED";
    FD1P3AX key_mem_14___i338 (.D(key_mem_0__127__N_6496[81]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [81])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i338.GSR = "ENABLED";
    FD1P3AX key_mem_14___i339 (.D(key_mem_0__127__N_6496[82]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [82])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i339.GSR = "ENABLED";
    FD1P3AX key_mem_14___i340 (.D(key_mem_0__127__N_6496[83]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [83])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i340.GSR = "ENABLED";
    FD1P3AX key_mem_14___i341 (.D(key_mem_0__127__N_6496[84]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [84])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i341.GSR = "ENABLED";
    FD1P3AX key_mem_14___i342 (.D(key_mem_0__127__N_6496[85]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [85])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i342.GSR = "ENABLED";
    FD1P3AX key_mem_14___i343 (.D(key_mem_0__127__N_6496[86]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [86])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i343.GSR = "ENABLED";
    FD1P3AX key_mem_14___i344 (.D(key_mem_0__127__N_6496[87]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [87])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i344.GSR = "ENABLED";
    FD1P3AX key_mem_14___i345 (.D(key_mem_0__127__N_6496[88]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [88])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i345.GSR = "ENABLED";
    FD1P3AX key_mem_14___i346 (.D(key_mem_0__127__N_6496[89]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [89])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i346.GSR = "ENABLED";
    FD1P3AX key_mem_14___i347 (.D(key_mem_0__127__N_6496[90]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [90])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i347.GSR = "ENABLED";
    FD1P3AX key_mem_14___i348 (.D(key_mem_0__127__N_6496[91]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [91])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i348.GSR = "ENABLED";
    FD1P3AX key_mem_14___i349 (.D(key_mem_0__127__N_6496[92]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [92])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i349.GSR = "ENABLED";
    FD1P3AX key_mem_14___i350 (.D(key_mem_0__127__N_6496[93]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(\key_mem[12] [93])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i350.GSR = "ENABLED";
    FD1P3AX key_mem_14___i351 (.D(key_mem_0__127__N_6496[94]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[12] [94])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i351.GSR = "ENABLED";
    FD1P3AX key_mem_14___i352 (.D(key_mem_0__127__N_6496[95]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[12] [95])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i352.GSR = "ENABLED";
    FD1P3AX key_mem_14___i353 (.D(key_mem_0__127__N_6496[96]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[12] [96])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i353.GSR = "ENABLED";
    FD1P3AX key_mem_14___i354 (.D(key_mem_0__127__N_6496[97]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[12] [97])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i354.GSR = "ENABLED";
    FD1P3AX key_mem_14___i355 (.D(key_mem_0__127__N_6496[98]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[12] [98])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i355.GSR = "ENABLED";
    FD1P3AX key_mem_14___i356 (.D(key_mem_0__127__N_6496[99]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[12] [99])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i356.GSR = "ENABLED";
    FD1P3AX key_mem_14___i357 (.D(key_mem_0__127__N_6496[100]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[12] [100])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i357.GSR = "ENABLED";
    FD1P3AX key_mem_14___i358 (.D(key_mem_0__127__N_6496[101]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[12] [101])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i358.GSR = "ENABLED";
    FD1P3AX key_mem_14___i359 (.D(key_mem_0__127__N_6496[102]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[12] [102])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i359.GSR = "ENABLED";
    FD1P3AX key_mem_14___i360 (.D(key_mem_0__127__N_6496[103]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[12] [103])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i360.GSR = "ENABLED";
    FD1P3AX key_mem_14___i361 (.D(key_mem_0__127__N_6496[104]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[12] [104])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i361.GSR = "ENABLED";
    FD1P3AX key_mem_14___i362 (.D(key_mem_0__127__N_6496[105]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[12] [105])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i362.GSR = "ENABLED";
    FD1P3AX key_mem_14___i363 (.D(key_mem_0__127__N_6496[106]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[12] [106])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i363.GSR = "ENABLED";
    FD1P3AX key_mem_14___i364 (.D(key_mem_0__127__N_6496[107]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[12] [107])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i364.GSR = "ENABLED";
    FD1P3AX key_mem_14___i365 (.D(key_mem_0__127__N_6496[108]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[12] [108])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i365.GSR = "ENABLED";
    FD1P3AX key_mem_14___i366 (.D(key_mem_0__127__N_6496[109]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[12] [109])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i366.GSR = "ENABLED";
    FD1P3AX key_mem_14___i367 (.D(key_mem_0__127__N_6496[110]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[12] [110])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i367.GSR = "ENABLED";
    FD1P3AX key_mem_14___i368 (.D(key_mem_0__127__N_6496[111]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[12] [111])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i368.GSR = "ENABLED";
    FD1P3AX key_mem_14___i369 (.D(key_mem_0__127__N_6496[112]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[12] [112])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i369.GSR = "ENABLED";
    FD1P3AX key_mem_14___i370 (.D(key_mem_0__127__N_6496[113]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[12] [113])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i370.GSR = "ENABLED";
    FD1P3AX key_mem_14___i371 (.D(key_mem_0__127__N_6496[114]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[12] [114])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i371.GSR = "ENABLED";
    FD1P3AX key_mem_14___i372 (.D(key_mem_0__127__N_6496[115]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[12] [115])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i372.GSR = "ENABLED";
    FD1P3AX key_mem_14___i373 (.D(key_mem_0__127__N_6496[116]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[12] [116])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i373.GSR = "ENABLED";
    FD1P3AX key_mem_14___i374 (.D(key_mem_0__127__N_6496[117]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[12] [117])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i374.GSR = "ENABLED";
    FD1P3AX key_mem_14___i375 (.D(key_mem_0__127__N_6496[118]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[12] [118])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i375.GSR = "ENABLED";
    FD1P3AX key_mem_14___i376 (.D(key_mem_0__127__N_6496[119]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[12] [119])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i376.GSR = "ENABLED";
    FD1P3AX key_mem_14___i377 (.D(key_mem_0__127__N_6496[120]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[12] [120])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i377.GSR = "ENABLED";
    FD1P3AX key_mem_14___i378 (.D(key_mem_0__127__N_6496[121]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[12] [121])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i378.GSR = "ENABLED";
    FD1P3AX key_mem_14___i379 (.D(key_mem_0__127__N_6496[122]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[12] [122])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i379.GSR = "ENABLED";
    FD1P3AX key_mem_14___i380 (.D(key_mem_0__127__N_6496[123]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[12] [123])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i380.GSR = "ENABLED";
    FD1P3AX key_mem_14___i381 (.D(key_mem_0__127__N_6496[124]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[12] [124])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i381.GSR = "ENABLED";
    FD1P3AX key_mem_14___i382 (.D(key_mem_0__127__N_6496[125]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[12] [125])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i382.GSR = "ENABLED";
    FD1P3AX key_mem_14___i383 (.D(key_mem_0__127__N_6496[126]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[12] [126])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i383.GSR = "ENABLED";
    FD1P3AX key_mem_14___i384 (.D(key_mem_0__127__N_6496[127]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[12] [127])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i384.GSR = "ENABLED";
    FD1P3AX key_mem_14___i385 (.D(key_mem_0__127__N_6368[0]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[11] [0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i385.GSR = "ENABLED";
    FD1P3AX key_mem_14___i386 (.D(key_mem_0__127__N_6368[1]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[11] [1])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i386.GSR = "ENABLED";
    FD1P3AX key_mem_14___i387 (.D(key_mem_0__127__N_6368[2]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[11] [2])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i387.GSR = "ENABLED";
    FD1P3AX key_mem_14___i388 (.D(key_mem_0__127__N_6368[3]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[11] [3])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i388.GSR = "ENABLED";
    FD1P3AX key_mem_14___i389 (.D(key_mem_0__127__N_6368[4]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[11] [4])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i389.GSR = "ENABLED";
    FD1P3AX key_mem_14___i390 (.D(key_mem_0__127__N_6368[5]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[11] [5])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i390.GSR = "ENABLED";
    FD1P3AX key_mem_14___i391 (.D(key_mem_0__127__N_6368[6]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[11] [6])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i391.GSR = "ENABLED";
    FD1P3AX key_mem_14___i392 (.D(key_mem_0__127__N_6368[7]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[11] [7])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i392.GSR = "ENABLED";
    FD1P3AX key_mem_14___i393 (.D(key_mem_0__127__N_6368[8]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[11] [8])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i393.GSR = "ENABLED";
    FD1P3AX key_mem_14___i394 (.D(key_mem_0__127__N_6368[9]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[11] [9])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i394.GSR = "ENABLED";
    FD1P3AX key_mem_14___i395 (.D(key_mem_0__127__N_6368[10]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[11] [10])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i395.GSR = "ENABLED";
    FD1P3AX key_mem_14___i396 (.D(key_mem_0__127__N_6368[11]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[11] [11])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i396.GSR = "ENABLED";
    FD1P3AX key_mem_14___i397 (.D(key_mem_0__127__N_6368[12]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[11] [12])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i397.GSR = "ENABLED";
    FD1P3AX key_mem_14___i398 (.D(key_mem_0__127__N_6368[13]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[11] [13])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i398.GSR = "ENABLED";
    FD1P3AX key_mem_14___i399 (.D(key_mem_0__127__N_6368[14]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[11] [14])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i399.GSR = "ENABLED";
    FD1P3AX key_mem_14___i400 (.D(key_mem_0__127__N_6368[15]), .SP(clk_c_enable_786), 
            .CK(clk_c), .Q(\key_mem[11] [15])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i400.GSR = "ENABLED";
    FD1P3AX key_mem_14___i401 (.D(key_mem_0__127__N_6368[16]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [16])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i401.GSR = "ENABLED";
    FD1P3AX key_mem_14___i402 (.D(key_mem_0__127__N_6368[17]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [17])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i402.GSR = "ENABLED";
    FD1P3AX key_mem_14___i403 (.D(key_mem_0__127__N_6368[18]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [18])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i403.GSR = "ENABLED";
    FD1P3AX key_mem_14___i404 (.D(key_mem_0__127__N_6368[19]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [19])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i404.GSR = "ENABLED";
    FD1P3AX key_mem_14___i405 (.D(key_mem_0__127__N_6368[20]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [20])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i405.GSR = "ENABLED";
    FD1P3AX key_mem_14___i406 (.D(key_mem_0__127__N_6368[21]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [21])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i406.GSR = "ENABLED";
    FD1P3AX key_mem_14___i407 (.D(key_mem_0__127__N_6368[22]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [22])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i407.GSR = "ENABLED";
    FD1P3AX key_mem_14___i408 (.D(key_mem_0__127__N_6368[23]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [23])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i408.GSR = "ENABLED";
    FD1P3AX key_mem_14___i409 (.D(key_mem_0__127__N_6368[24]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [24])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i409.GSR = "ENABLED";
    FD1P3AX key_mem_14___i410 (.D(key_mem_0__127__N_6368[25]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [25])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i410.GSR = "ENABLED";
    FD1P3AX key_mem_14___i411 (.D(key_mem_0__127__N_6368[26]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [26])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i411.GSR = "ENABLED";
    FD1P3AX key_mem_14___i412 (.D(key_mem_0__127__N_6368[27]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [27])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i412.GSR = "ENABLED";
    FD1P3AX key_mem_14___i413 (.D(key_mem_0__127__N_6368[28]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [28])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i413.GSR = "ENABLED";
    FD1P3AX key_mem_14___i414 (.D(key_mem_0__127__N_6368[29]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [29])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i414.GSR = "ENABLED";
    FD1P3AX key_mem_14___i415 (.D(key_mem_0__127__N_6368[30]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [30])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i415.GSR = "ENABLED";
    FD1P3AX key_mem_14___i416 (.D(key_mem_0__127__N_6368[31]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [31])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i416.GSR = "ENABLED";
    FD1P3AX key_mem_14___i417 (.D(key_mem_0__127__N_6368[32]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [32])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i417.GSR = "ENABLED";
    FD1P3AX key_mem_14___i418 (.D(key_mem_0__127__N_6368[33]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [33])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i418.GSR = "ENABLED";
    FD1P3AX key_mem_14___i419 (.D(key_mem_0__127__N_6368[34]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [34])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i419.GSR = "ENABLED";
    FD1P3AX key_mem_14___i420 (.D(key_mem_0__127__N_6368[35]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [35])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i420.GSR = "ENABLED";
    FD1P3AX key_mem_14___i421 (.D(key_mem_0__127__N_6368[36]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [36])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i421.GSR = "ENABLED";
    FD1P3AX key_mem_14___i422 (.D(key_mem_0__127__N_6368[37]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [37])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i422.GSR = "ENABLED";
    FD1P3AX key_mem_14___i423 (.D(key_mem_0__127__N_6368[38]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [38])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i423.GSR = "ENABLED";
    FD1P3AX key_mem_14___i424 (.D(key_mem_0__127__N_6368[39]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [39])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i424.GSR = "ENABLED";
    FD1P3AX key_mem_14___i425 (.D(key_mem_0__127__N_6368[40]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [40])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i425.GSR = "ENABLED";
    FD1P3AX key_mem_14___i426 (.D(key_mem_0__127__N_6368[41]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [41])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i426.GSR = "ENABLED";
    FD1P3AX key_mem_14___i427 (.D(key_mem_0__127__N_6368[42]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [42])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i427.GSR = "ENABLED";
    FD1P3AX key_mem_14___i428 (.D(key_mem_0__127__N_6368[43]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [43])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i428.GSR = "ENABLED";
    FD1P3AX key_mem_14___i429 (.D(key_mem_0__127__N_6368[44]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [44])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i429.GSR = "ENABLED";
    FD1P3AX key_mem_14___i430 (.D(key_mem_0__127__N_6368[45]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [45])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i430.GSR = "ENABLED";
    FD1P3AX key_mem_14___i431 (.D(key_mem_0__127__N_6368[46]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [46])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i431.GSR = "ENABLED";
    FD1P3AX key_mem_14___i432 (.D(key_mem_0__127__N_6368[47]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [47])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i432.GSR = "ENABLED";
    FD1P3AX key_mem_14___i433 (.D(key_mem_0__127__N_6368[48]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [48])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i433.GSR = "ENABLED";
    FD1P3AX key_mem_14___i434 (.D(key_mem_0__127__N_6368[49]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [49])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i434.GSR = "ENABLED";
    FD1P3AX key_mem_14___i435 (.D(key_mem_0__127__N_6368[50]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [50])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i435.GSR = "ENABLED";
    FD1P3AX key_mem_14___i436 (.D(key_mem_0__127__N_6368[51]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [51])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i436.GSR = "ENABLED";
    FD1P3AX key_mem_14___i437 (.D(key_mem_0__127__N_6368[52]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [52])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i437.GSR = "ENABLED";
    FD1P3AX key_mem_14___i438 (.D(key_mem_0__127__N_6368[53]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [53])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i438.GSR = "ENABLED";
    FD1P3AX key_mem_14___i439 (.D(key_mem_0__127__N_6368[54]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [54])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i439.GSR = "ENABLED";
    FD1P3AX key_mem_14___i440 (.D(key_mem_0__127__N_6368[55]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [55])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i440.GSR = "ENABLED";
    FD1P3AX key_mem_14___i441 (.D(key_mem_0__127__N_6368[56]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [56])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i441.GSR = "ENABLED";
    FD1P3AX key_mem_14___i442 (.D(key_mem_0__127__N_6368[57]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [57])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i442.GSR = "ENABLED";
    FD1P3AX key_mem_14___i443 (.D(key_mem_0__127__N_6368[58]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [58])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i443.GSR = "ENABLED";
    FD1P3AX key_mem_14___i444 (.D(key_mem_0__127__N_6368[59]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [59])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i444.GSR = "ENABLED";
    FD1P3AX key_mem_14___i445 (.D(key_mem_0__127__N_6368[60]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [60])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i445.GSR = "ENABLED";
    FD1P3AX key_mem_14___i446 (.D(key_mem_0__127__N_6368[61]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [61])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i446.GSR = "ENABLED";
    FD1P3AX key_mem_14___i447 (.D(key_mem_0__127__N_6368[62]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [62])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i447.GSR = "ENABLED";
    FD1P3AX key_mem_14___i448 (.D(key_mem_0__127__N_6368[63]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [63])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i448.GSR = "ENABLED";
    FD1P3AX key_mem_14___i449 (.D(key_mem_0__127__N_6368[64]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [64])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i449.GSR = "ENABLED";
    FD1P3AX key_mem_14___i450 (.D(key_mem_0__127__N_6368[65]), .SP(clk_c_enable_836), 
            .CK(clk_c), .Q(\key_mem[11] [65])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i450.GSR = "ENABLED";
    FD1P3AX key_mem_14___i451 (.D(key_mem_0__127__N_6368[66]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [66])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i451.GSR = "ENABLED";
    FD1P3AX key_mem_14___i452 (.D(key_mem_0__127__N_6368[67]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [67])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i452.GSR = "ENABLED";
    FD1P3AX key_mem_14___i453 (.D(key_mem_0__127__N_6368[68]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [68])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i453.GSR = "ENABLED";
    FD1P3AX key_mem_14___i454 (.D(key_mem_0__127__N_6368[69]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [69])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i454.GSR = "ENABLED";
    FD1P3AX key_mem_14___i455 (.D(key_mem_0__127__N_6368[70]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [70])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i455.GSR = "ENABLED";
    FD1P3AX key_mem_14___i456 (.D(key_mem_0__127__N_6368[71]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [71])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i456.GSR = "ENABLED";
    FD1P3AX key_mem_14___i457 (.D(key_mem_0__127__N_6368[72]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [72])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i457.GSR = "ENABLED";
    FD1P3AX key_mem_14___i458 (.D(key_mem_0__127__N_6368[73]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [73])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i458.GSR = "ENABLED";
    FD1P3AX key_mem_14___i459 (.D(key_mem_0__127__N_6368[74]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [74])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i459.GSR = "ENABLED";
    FD1P3AX key_mem_14___i460 (.D(key_mem_0__127__N_6368[75]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [75])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i460.GSR = "ENABLED";
    FD1P3AX key_mem_14___i461 (.D(key_mem_0__127__N_6368[76]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [76])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i461.GSR = "ENABLED";
    FD1P3AX key_mem_14___i462 (.D(key_mem_0__127__N_6368[77]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [77])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i462.GSR = "ENABLED";
    FD1P3AX key_mem_14___i463 (.D(key_mem_0__127__N_6368[78]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [78])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i463.GSR = "ENABLED";
    FD1P3AX key_mem_14___i464 (.D(key_mem_0__127__N_6368[79]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [79])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i464.GSR = "ENABLED";
    FD1P3AX key_mem_14___i465 (.D(key_mem_0__127__N_6368[80]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [80])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i465.GSR = "ENABLED";
    FD1P3AX key_mem_14___i466 (.D(key_mem_0__127__N_6368[81]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [81])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i466.GSR = "ENABLED";
    FD1P3AX key_mem_14___i467 (.D(key_mem_0__127__N_6368[82]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [82])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i467.GSR = "ENABLED";
    FD1P3AX key_mem_14___i468 (.D(key_mem_0__127__N_6368[83]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [83])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i468.GSR = "ENABLED";
    FD1P3AX key_mem_14___i469 (.D(key_mem_0__127__N_6368[84]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [84])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i469.GSR = "ENABLED";
    FD1P3AX key_mem_14___i470 (.D(key_mem_0__127__N_6368[85]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [85])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i470.GSR = "ENABLED";
    FD1P3AX key_mem_14___i471 (.D(key_mem_0__127__N_6368[86]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [86])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i471.GSR = "ENABLED";
    FD1P3AX key_mem_14___i472 (.D(key_mem_0__127__N_6368[87]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [87])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i472.GSR = "ENABLED";
    FD1P3AX key_mem_14___i473 (.D(key_mem_0__127__N_6368[88]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [88])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i473.GSR = "ENABLED";
    FD1P3AX key_mem_14___i474 (.D(key_mem_0__127__N_6368[89]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [89])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i474.GSR = "ENABLED";
    FD1P3AX key_mem_14___i475 (.D(key_mem_0__127__N_6368[90]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [90])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i475.GSR = "ENABLED";
    FD1P3AX key_mem_14___i476 (.D(key_mem_0__127__N_6368[91]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [91])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i476.GSR = "ENABLED";
    FD1P3AX key_mem_14___i477 (.D(key_mem_0__127__N_6368[92]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [92])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i477.GSR = "ENABLED";
    FD1P3AX key_mem_14___i478 (.D(key_mem_0__127__N_6368[93]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [93])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i478.GSR = "ENABLED";
    FD1P3AX key_mem_14___i479 (.D(key_mem_0__127__N_6368[94]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [94])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i479.GSR = "ENABLED";
    FD1P3AX key_mem_14___i480 (.D(key_mem_0__127__N_6368[95]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [95])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i480.GSR = "ENABLED";
    FD1P3AX key_mem_14___i481 (.D(key_mem_0__127__N_6368[96]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [96])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i481.GSR = "ENABLED";
    FD1P3AX key_mem_14___i482 (.D(key_mem_0__127__N_6368[97]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [97])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i482.GSR = "ENABLED";
    FD1P3AX key_mem_14___i483 (.D(key_mem_0__127__N_6368[98]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [98])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i483.GSR = "ENABLED";
    FD1P3AX key_mem_14___i484 (.D(key_mem_0__127__N_6368[99]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [99])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i484.GSR = "ENABLED";
    FD1P3AX key_mem_14___i485 (.D(key_mem_0__127__N_6368[100]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [100])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i485.GSR = "ENABLED";
    FD1P3AX key_mem_14___i486 (.D(key_mem_0__127__N_6368[101]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [101])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i486.GSR = "ENABLED";
    FD1P3AX key_mem_14___i487 (.D(key_mem_0__127__N_6368[102]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [102])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i487.GSR = "ENABLED";
    FD1P3AX key_mem_14___i488 (.D(key_mem_0__127__N_6368[103]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [103])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i488.GSR = "ENABLED";
    FD1P3AX key_mem_14___i489 (.D(key_mem_0__127__N_6368[104]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [104])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i489.GSR = "ENABLED";
    FD1P3AX key_mem_14___i490 (.D(key_mem_0__127__N_6368[105]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [105])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i490.GSR = "ENABLED";
    FD1P3AX key_mem_14___i491 (.D(key_mem_0__127__N_6368[106]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [106])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i491.GSR = "ENABLED";
    FD1P3AX key_mem_14___i492 (.D(key_mem_0__127__N_6368[107]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [107])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i492.GSR = "ENABLED";
    FD1P3AX key_mem_14___i493 (.D(key_mem_0__127__N_6368[108]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [108])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i493.GSR = "ENABLED";
    FD1P3AX key_mem_14___i494 (.D(key_mem_0__127__N_6368[109]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [109])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i494.GSR = "ENABLED";
    FD1P3AX key_mem_14___i495 (.D(key_mem_0__127__N_6368[110]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [110])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i495.GSR = "ENABLED";
    FD1P3AX key_mem_14___i496 (.D(key_mem_0__127__N_6368[111]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [111])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i496.GSR = "ENABLED";
    FD1P3AX key_mem_14___i497 (.D(key_mem_0__127__N_6368[112]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [112])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i497.GSR = "ENABLED";
    FD1P3AX key_mem_14___i498 (.D(key_mem_0__127__N_6368[113]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [113])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i498.GSR = "ENABLED";
    FD1P3AX key_mem_14___i499 (.D(key_mem_0__127__N_6368[114]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [114])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i499.GSR = "ENABLED";
    FD1P3AX key_mem_14___i500 (.D(key_mem_0__127__N_6368[115]), .SP(clk_c_enable_886), 
            .CK(clk_c), .Q(\key_mem[11] [115])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i500.GSR = "ENABLED";
    FD1P3AX key_mem_14___i501 (.D(key_mem_0__127__N_6368[116]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[11] [116])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i501.GSR = "ENABLED";
    FD1P3AX key_mem_14___i502 (.D(key_mem_0__127__N_6368[117]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[11] [117])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i502.GSR = "ENABLED";
    FD1P3AX key_mem_14___i503 (.D(key_mem_0__127__N_6368[118]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[11] [118])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i503.GSR = "ENABLED";
    FD1P3AX key_mem_14___i504 (.D(key_mem_0__127__N_6368[119]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[11] [119])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i504.GSR = "ENABLED";
    FD1P3AX key_mem_14___i505 (.D(key_mem_0__127__N_6368[120]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[11] [120])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i505.GSR = "ENABLED";
    FD1P3AX key_mem_14___i506 (.D(key_mem_0__127__N_6368[121]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[11] [121])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i506.GSR = "ENABLED";
    FD1P3AX key_mem_14___i507 (.D(key_mem_0__127__N_6368[122]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[11] [122])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i507.GSR = "ENABLED";
    FD1P3AX key_mem_14___i508 (.D(key_mem_0__127__N_6368[123]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[11] [123])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i508.GSR = "ENABLED";
    FD1P3AX key_mem_14___i509 (.D(key_mem_0__127__N_6368[124]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[11] [124])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i509.GSR = "ENABLED";
    FD1P3AX key_mem_14___i510 (.D(key_mem_0__127__N_6368[125]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[11] [125])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i510.GSR = "ENABLED";
    FD1P3AX key_mem_14___i511 (.D(key_mem_0__127__N_6368[126]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[11] [126])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i511.GSR = "ENABLED";
    FD1P3AX key_mem_14___i512 (.D(key_mem_0__127__N_6368[127]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[11] [127])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i512.GSR = "ENABLED";
    FD1P3AX key_mem_14___i513 (.D(key_mem_0__127__N_6240[0]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[10] [0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i513.GSR = "ENABLED";
    FD1P3AX key_mem_14___i514 (.D(key_mem_0__127__N_6240[1]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[10] [1])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i514.GSR = "ENABLED";
    FD1P3AX key_mem_14___i515 (.D(key_mem_0__127__N_6240[2]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[10] [2])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i515.GSR = "ENABLED";
    FD1P3AX key_mem_14___i516 (.D(key_mem_0__127__N_6240[3]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[10] [3])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i516.GSR = "ENABLED";
    FD1P3AX key_mem_14___i517 (.D(key_mem_0__127__N_6240[4]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[10] [4])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i517.GSR = "ENABLED";
    FD1P3AX key_mem_14___i518 (.D(key_mem_0__127__N_6240[5]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[10] [5])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i518.GSR = "ENABLED";
    FD1P3AX key_mem_14___i519 (.D(key_mem_0__127__N_6240[6]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[10] [6])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i519.GSR = "ENABLED";
    FD1P3AX key_mem_14___i520 (.D(key_mem_0__127__N_6240[7]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[10] [7])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i520.GSR = "ENABLED";
    FD1P3AX key_mem_14___i521 (.D(key_mem_0__127__N_6240[8]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[10] [8])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i521.GSR = "ENABLED";
    FD1P3AX key_mem_14___i522 (.D(key_mem_0__127__N_6240[9]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[10] [9])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i522.GSR = "ENABLED";
    FD1P3AX key_mem_14___i523 (.D(key_mem_0__127__N_6240[10]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[10] [10])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i523.GSR = "ENABLED";
    FD1P3AX key_mem_14___i524 (.D(key_mem_0__127__N_6240[11]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[10] [11])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i524.GSR = "ENABLED";
    FD1P3AX key_mem_14___i525 (.D(key_mem_0__127__N_6240[12]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[10] [12])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i525.GSR = "ENABLED";
    FD1P3AX key_mem_14___i526 (.D(key_mem_0__127__N_6240[13]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[10] [13])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i526.GSR = "ENABLED";
    FD1P3AX key_mem_14___i527 (.D(key_mem_0__127__N_6240[14]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[10] [14])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i527.GSR = "ENABLED";
    FD1P3AX key_mem_14___i528 (.D(key_mem_0__127__N_6240[15]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[10] [15])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i528.GSR = "ENABLED";
    FD1P3AX key_mem_14___i529 (.D(key_mem_0__127__N_6240[16]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[10] [16])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i529.GSR = "ENABLED";
    FD1P3AX key_mem_14___i530 (.D(key_mem_0__127__N_6240[17]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[10] [17])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i530.GSR = "ENABLED";
    FD1P3AX key_mem_14___i531 (.D(key_mem_0__127__N_6240[18]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[10] [18])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i531.GSR = "ENABLED";
    FD1P3AX key_mem_14___i532 (.D(key_mem_0__127__N_6240[19]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[10] [19])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i532.GSR = "ENABLED";
    FD1P3AX key_mem_14___i533 (.D(key_mem_0__127__N_6240[20]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[10] [20])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i533.GSR = "ENABLED";
    FD1P3AX key_mem_14___i534 (.D(key_mem_0__127__N_6240[21]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[10] [21])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i534.GSR = "ENABLED";
    FD1P3AX key_mem_14___i535 (.D(key_mem_0__127__N_6240[22]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[10] [22])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i535.GSR = "ENABLED";
    FD1P3AX key_mem_14___i536 (.D(key_mem_0__127__N_6240[23]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[10] [23])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i536.GSR = "ENABLED";
    FD1P3AX key_mem_14___i537 (.D(key_mem_0__127__N_6240[24]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[10] [24])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i537.GSR = "ENABLED";
    FD1P3AX key_mem_14___i538 (.D(key_mem_0__127__N_6240[25]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[10] [25])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i538.GSR = "ENABLED";
    FD1P3AX key_mem_14___i539 (.D(key_mem_0__127__N_6240[26]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[10] [26])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i539.GSR = "ENABLED";
    FD1P3AX key_mem_14___i540 (.D(key_mem_0__127__N_6240[27]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[10] [27])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i540.GSR = "ENABLED";
    FD1P3AX key_mem_14___i541 (.D(key_mem_0__127__N_6240[28]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[10] [28])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i541.GSR = "ENABLED";
    FD1P3AX key_mem_14___i542 (.D(key_mem_0__127__N_6240[29]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[10] [29])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i542.GSR = "ENABLED";
    FD1P3AX key_mem_14___i543 (.D(key_mem_0__127__N_6240[30]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[10] [30])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i543.GSR = "ENABLED";
    FD1P3AX key_mem_14___i544 (.D(key_mem_0__127__N_6240[31]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[10] [31])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i544.GSR = "ENABLED";
    FD1P3AX key_mem_14___i545 (.D(key_mem_0__127__N_6240[32]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[10] [32])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i545.GSR = "ENABLED";
    FD1P3AX key_mem_14___i546 (.D(key_mem_0__127__N_6240[33]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[10] [33])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i546.GSR = "ENABLED";
    FD1P3AX key_mem_14___i547 (.D(key_mem_0__127__N_6240[34]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[10] [34])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i547.GSR = "ENABLED";
    FD1P3AX key_mem_14___i548 (.D(key_mem_0__127__N_6240[35]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[10] [35])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i548.GSR = "ENABLED";
    FD1P3AX key_mem_14___i549 (.D(key_mem_0__127__N_6240[36]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[10] [36])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i549.GSR = "ENABLED";
    FD1P3AX key_mem_14___i550 (.D(key_mem_0__127__N_6240[37]), .SP(clk_c_enable_936), 
            .CK(clk_c), .Q(\key_mem[10] [37])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i550.GSR = "ENABLED";
    FD1P3AX key_mem_14___i551 (.D(key_mem_0__127__N_6240[38]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [38])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i551.GSR = "ENABLED";
    FD1P3AX key_mem_14___i552 (.D(key_mem_0__127__N_6240[39]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [39])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i552.GSR = "ENABLED";
    FD1P3AX key_mem_14___i553 (.D(key_mem_0__127__N_6240[40]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [40])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i553.GSR = "ENABLED";
    FD1P3AX key_mem_14___i554 (.D(key_mem_0__127__N_6240[41]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [41])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i554.GSR = "ENABLED";
    FD1P3AX key_mem_14___i555 (.D(key_mem_0__127__N_6240[42]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [42])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i555.GSR = "ENABLED";
    FD1P3AX key_mem_14___i556 (.D(key_mem_0__127__N_6240[43]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [43])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i556.GSR = "ENABLED";
    FD1P3AX key_mem_14___i557 (.D(key_mem_0__127__N_6240[44]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [44])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i557.GSR = "ENABLED";
    FD1P3AX key_mem_14___i558 (.D(key_mem_0__127__N_6240[45]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [45])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i558.GSR = "ENABLED";
    FD1P3AX key_mem_14___i559 (.D(key_mem_0__127__N_6240[46]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [46])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i559.GSR = "ENABLED";
    FD1P3AX key_mem_14___i560 (.D(key_mem_0__127__N_6240[47]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [47])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i560.GSR = "ENABLED";
    FD1P3AX key_mem_14___i561 (.D(key_mem_0__127__N_6240[48]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [48])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i561.GSR = "ENABLED";
    FD1P3AX key_mem_14___i562 (.D(key_mem_0__127__N_6240[49]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [49])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i562.GSR = "ENABLED";
    FD1P3AX key_mem_14___i563 (.D(key_mem_0__127__N_6240[50]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [50])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i563.GSR = "ENABLED";
    FD1P3AX key_mem_14___i564 (.D(key_mem_0__127__N_6240[51]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [51])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i564.GSR = "ENABLED";
    FD1P3AX key_mem_14___i565 (.D(key_mem_0__127__N_6240[52]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [52])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i565.GSR = "ENABLED";
    FD1P3AX key_mem_14___i566 (.D(key_mem_0__127__N_6240[53]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [53])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i566.GSR = "ENABLED";
    FD1P3AX key_mem_14___i567 (.D(key_mem_0__127__N_6240[54]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [54])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i567.GSR = "ENABLED";
    FD1P3AX key_mem_14___i568 (.D(key_mem_0__127__N_6240[55]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [55])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i568.GSR = "ENABLED";
    FD1P3AX key_mem_14___i569 (.D(key_mem_0__127__N_6240[56]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [56])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i569.GSR = "ENABLED";
    FD1P3AX key_mem_14___i570 (.D(key_mem_0__127__N_6240[57]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [57])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i570.GSR = "ENABLED";
    FD1P3AX key_mem_14___i571 (.D(key_mem_0__127__N_6240[58]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [58])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i571.GSR = "ENABLED";
    FD1P3AX key_mem_14___i572 (.D(key_mem_0__127__N_6240[59]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [59])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i572.GSR = "ENABLED";
    FD1P3AX key_mem_14___i573 (.D(key_mem_0__127__N_6240[60]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [60])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i573.GSR = "ENABLED";
    FD1P3AX key_mem_14___i574 (.D(key_mem_0__127__N_6240[61]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [61])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i574.GSR = "ENABLED";
    FD1P3AX key_mem_14___i575 (.D(key_mem_0__127__N_6240[62]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [62])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i575.GSR = "ENABLED";
    FD1P3AX key_mem_14___i576 (.D(key_mem_0__127__N_6240[63]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [63])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i576.GSR = "ENABLED";
    FD1P3AX key_mem_14___i577 (.D(key_mem_0__127__N_6240[64]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [64])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i577.GSR = "ENABLED";
    FD1P3AX key_mem_14___i578 (.D(key_mem_0__127__N_6240[65]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [65])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i578.GSR = "ENABLED";
    FD1P3AX key_mem_14___i579 (.D(key_mem_0__127__N_6240[66]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [66])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i579.GSR = "ENABLED";
    FD1P3AX key_mem_14___i580 (.D(key_mem_0__127__N_6240[67]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [67])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i580.GSR = "ENABLED";
    FD1P3AX key_mem_14___i581 (.D(key_mem_0__127__N_6240[68]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [68])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i581.GSR = "ENABLED";
    FD1P3AX key_mem_14___i582 (.D(key_mem_0__127__N_6240[69]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [69])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i582.GSR = "ENABLED";
    FD1P3AX key_mem_14___i583 (.D(key_mem_0__127__N_6240[70]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [70])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i583.GSR = "ENABLED";
    FD1P3AX key_mem_14___i584 (.D(key_mem_0__127__N_6240[71]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [71])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i584.GSR = "ENABLED";
    FD1P3AX key_mem_14___i585 (.D(key_mem_0__127__N_6240[72]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [72])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i585.GSR = "ENABLED";
    FD1P3AX key_mem_14___i586 (.D(key_mem_0__127__N_6240[73]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [73])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i586.GSR = "ENABLED";
    FD1P3AX key_mem_14___i587 (.D(key_mem_0__127__N_6240[74]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [74])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i587.GSR = "ENABLED";
    FD1P3AX key_mem_14___i588 (.D(key_mem_0__127__N_6240[75]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [75])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i588.GSR = "ENABLED";
    FD1P3AX key_mem_14___i589 (.D(key_mem_0__127__N_6240[76]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [76])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i589.GSR = "ENABLED";
    FD1P3AX key_mem_14___i590 (.D(key_mem_0__127__N_6240[77]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [77])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i590.GSR = "ENABLED";
    FD1P3AX key_mem_14___i591 (.D(key_mem_0__127__N_6240[78]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [78])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i591.GSR = "ENABLED";
    FD1P3AX key_mem_14___i592 (.D(key_mem_0__127__N_6240[79]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [79])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i592.GSR = "ENABLED";
    FD1P3AX key_mem_14___i593 (.D(key_mem_0__127__N_6240[80]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [80])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i593.GSR = "ENABLED";
    FD1P3AX key_mem_14___i594 (.D(key_mem_0__127__N_6240[81]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [81])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i594.GSR = "ENABLED";
    FD1P3AX key_mem_14___i595 (.D(key_mem_0__127__N_6240[82]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [82])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i595.GSR = "ENABLED";
    FD1P3AX key_mem_14___i596 (.D(key_mem_0__127__N_6240[83]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [83])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i596.GSR = "ENABLED";
    FD1P3AX key_mem_14___i597 (.D(key_mem_0__127__N_6240[84]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [84])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i597.GSR = "ENABLED";
    FD1P3AX key_mem_14___i598 (.D(key_mem_0__127__N_6240[85]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [85])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i598.GSR = "ENABLED";
    FD1P3AX key_mem_14___i599 (.D(key_mem_0__127__N_6240[86]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [86])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i599.GSR = "ENABLED";
    FD1P3AX key_mem_14___i600 (.D(key_mem_0__127__N_6240[87]), .SP(clk_c_enable_986), 
            .CK(clk_c), .Q(\key_mem[10] [87])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i600.GSR = "ENABLED";
    FD1P3AX key_mem_14___i601 (.D(key_mem_0__127__N_6240[88]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[10] [88])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i601.GSR = "ENABLED";
    FD1P3AX key_mem_14___i602 (.D(key_mem_0__127__N_6240[89]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[10] [89])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i602.GSR = "ENABLED";
    FD1P3AX key_mem_14___i603 (.D(key_mem_0__127__N_6240[90]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[10] [90])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i603.GSR = "ENABLED";
    FD1P3AX key_mem_14___i604 (.D(key_mem_0__127__N_6240[91]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[10] [91])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i604.GSR = "ENABLED";
    FD1P3AX key_mem_14___i605 (.D(key_mem_0__127__N_6240[92]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[10] [92])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i605.GSR = "ENABLED";
    FD1P3AX key_mem_14___i606 (.D(key_mem_0__127__N_6240[93]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[10] [93])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i606.GSR = "ENABLED";
    FD1P3AX key_mem_14___i607 (.D(key_mem_0__127__N_6240[94]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[10] [94])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i607.GSR = "ENABLED";
    FD1P3AX key_mem_14___i608 (.D(key_mem_0__127__N_6240[95]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[10] [95])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i608.GSR = "ENABLED";
    FD1P3AX key_mem_14___i609 (.D(key_mem_0__127__N_6240[96]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[10] [96])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i609.GSR = "ENABLED";
    FD1P3AX key_mem_14___i610 (.D(key_mem_0__127__N_6240[97]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[10] [97])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i610.GSR = "ENABLED";
    FD1P3AX key_mem_14___i611 (.D(key_mem_0__127__N_6240[98]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[10] [98])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i611.GSR = "ENABLED";
    FD1P3AX key_mem_14___i612 (.D(key_mem_0__127__N_6240[99]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[10] [99])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i612.GSR = "ENABLED";
    FD1P3AX key_mem_14___i613 (.D(key_mem_0__127__N_6240[100]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[10] [100])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i613.GSR = "ENABLED";
    FD1P3AX key_mem_14___i614 (.D(key_mem_0__127__N_6240[101]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[10] [101])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i614.GSR = "ENABLED";
    FD1P3AX key_mem_14___i615 (.D(key_mem_0__127__N_6240[102]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[10] [102])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i615.GSR = "ENABLED";
    FD1P3AX key_mem_14___i616 (.D(key_mem_0__127__N_6240[103]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[10] [103])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i616.GSR = "ENABLED";
    FD1P3AX key_mem_14___i617 (.D(key_mem_0__127__N_6240[104]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[10] [104])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i617.GSR = "ENABLED";
    FD1P3AX key_mem_14___i618 (.D(key_mem_0__127__N_6240[105]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[10] [105])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i618.GSR = "ENABLED";
    FD1P3AX key_mem_14___i619 (.D(key_mem_0__127__N_6240[106]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[10] [106])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i619.GSR = "ENABLED";
    FD1P3AX key_mem_14___i620 (.D(key_mem_0__127__N_6240[107]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[10] [107])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i620.GSR = "ENABLED";
    FD1P3AX key_mem_14___i621 (.D(key_mem_0__127__N_6240[108]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[10] [108])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i621.GSR = "ENABLED";
    FD1P3AX key_mem_14___i622 (.D(key_mem_0__127__N_6240[109]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[10] [109])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i622.GSR = "ENABLED";
    FD1P3AX key_mem_14___i623 (.D(key_mem_0__127__N_6240[110]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[10] [110])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i623.GSR = "ENABLED";
    FD1P3AX key_mem_14___i624 (.D(key_mem_0__127__N_6240[111]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[10] [111])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i624.GSR = "ENABLED";
    FD1P3AX key_mem_14___i625 (.D(key_mem_0__127__N_6240[112]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[10] [112])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i625.GSR = "ENABLED";
    FD1P3AX key_mem_14___i626 (.D(key_mem_0__127__N_6240[113]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[10] [113])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i626.GSR = "ENABLED";
    FD1P3AX key_mem_14___i627 (.D(key_mem_0__127__N_6240[114]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[10] [114])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i627.GSR = "ENABLED";
    FD1P3AX key_mem_14___i628 (.D(key_mem_0__127__N_6240[115]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[10] [115])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i628.GSR = "ENABLED";
    FD1P3AX key_mem_14___i629 (.D(key_mem_0__127__N_6240[116]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[10] [116])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i629.GSR = "ENABLED";
    FD1P3AX key_mem_14___i630 (.D(key_mem_0__127__N_6240[117]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[10] [117])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i630.GSR = "ENABLED";
    FD1P3AX key_mem_14___i631 (.D(key_mem_0__127__N_6240[118]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[10] [118])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i631.GSR = "ENABLED";
    FD1P3AX key_mem_14___i632 (.D(key_mem_0__127__N_6240[119]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[10] [119])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i632.GSR = "ENABLED";
    FD1P3AX key_mem_14___i633 (.D(key_mem_0__127__N_6240[120]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[10] [120])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i633.GSR = "ENABLED";
    FD1P3AX key_mem_14___i634 (.D(key_mem_0__127__N_6240[121]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[10] [121])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i634.GSR = "ENABLED";
    FD1P3AX key_mem_14___i635 (.D(key_mem_0__127__N_6240[122]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[10] [122])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i635.GSR = "ENABLED";
    FD1P3AX key_mem_14___i636 (.D(key_mem_0__127__N_6240[123]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[10] [123])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i636.GSR = "ENABLED";
    FD1P3AX key_mem_14___i637 (.D(key_mem_0__127__N_6240[124]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[10] [124])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i637.GSR = "ENABLED";
    FD1P3AX key_mem_14___i638 (.D(key_mem_0__127__N_6240[125]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[10] [125])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i638.GSR = "ENABLED";
    FD1P3AX key_mem_14___i639 (.D(key_mem_0__127__N_6240[126]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[10] [126])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i639.GSR = "ENABLED";
    FD1P3AX key_mem_14___i640 (.D(key_mem_0__127__N_6240[127]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[10] [127])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i640.GSR = "ENABLED";
    FD1P3AX key_mem_14___i641 (.D(key_mem_0__127__N_6112[0]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[9] [0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i641.GSR = "ENABLED";
    FD1P3AX key_mem_14___i642 (.D(key_mem_0__127__N_6112[1]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[9] [1])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i642.GSR = "ENABLED";
    FD1P3AX key_mem_14___i643 (.D(key_mem_0__127__N_6112[2]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[9] [2])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i643.GSR = "ENABLED";
    FD1P3AX key_mem_14___i644 (.D(key_mem_0__127__N_6112[3]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[9] [3])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i644.GSR = "ENABLED";
    FD1P3AX key_mem_14___i645 (.D(key_mem_0__127__N_6112[4]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[9] [4])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i645.GSR = "ENABLED";
    FD1P3AX key_mem_14___i646 (.D(key_mem_0__127__N_6112[5]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[9] [5])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i646.GSR = "ENABLED";
    FD1P3AX key_mem_14___i647 (.D(key_mem_0__127__N_6112[6]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[9] [6])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i647.GSR = "ENABLED";
    FD1P3AX key_mem_14___i648 (.D(key_mem_0__127__N_6112[7]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[9] [7])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i648.GSR = "ENABLED";
    FD1P3AX key_mem_14___i649 (.D(key_mem_0__127__N_6112[8]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[9] [8])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i649.GSR = "ENABLED";
    FD1P3AX key_mem_14___i650 (.D(key_mem_0__127__N_6112[9]), .SP(clk_c_enable_1036), 
            .CK(clk_c), .Q(\key_mem[9] [9])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i650.GSR = "ENABLED";
    FD1P3AX key_mem_14___i651 (.D(key_mem_0__127__N_6112[10]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [10])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i651.GSR = "ENABLED";
    FD1P3AX key_mem_14___i652 (.D(key_mem_0__127__N_6112[11]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [11])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i652.GSR = "ENABLED";
    FD1P3AX key_mem_14___i653 (.D(key_mem_0__127__N_6112[12]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [12])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i653.GSR = "ENABLED";
    FD1P3AX key_mem_14___i654 (.D(key_mem_0__127__N_6112[13]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [13])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i654.GSR = "ENABLED";
    FD1P3AX key_mem_14___i655 (.D(key_mem_0__127__N_6112[14]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [14])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i655.GSR = "ENABLED";
    FD1P3AX key_mem_14___i656 (.D(key_mem_0__127__N_6112[15]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [15])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i656.GSR = "ENABLED";
    FD1P3AX key_mem_14___i657 (.D(key_mem_0__127__N_6112[16]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [16])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i657.GSR = "ENABLED";
    FD1P3AX key_mem_14___i658 (.D(key_mem_0__127__N_6112[17]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [17])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i658.GSR = "ENABLED";
    FD1P3AX key_mem_14___i659 (.D(key_mem_0__127__N_6112[18]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [18])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i659.GSR = "ENABLED";
    FD1P3AX key_mem_14___i660 (.D(key_mem_0__127__N_6112[19]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [19])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i660.GSR = "ENABLED";
    FD1P3AX key_mem_14___i661 (.D(key_mem_0__127__N_6112[20]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [20])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i661.GSR = "ENABLED";
    FD1P3AX key_mem_14___i662 (.D(key_mem_0__127__N_6112[21]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [21])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i662.GSR = "ENABLED";
    FD1P3AX key_mem_14___i663 (.D(key_mem_0__127__N_6112[22]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [22])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i663.GSR = "ENABLED";
    FD1P3AX key_mem_14___i664 (.D(key_mem_0__127__N_6112[23]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [23])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i664.GSR = "ENABLED";
    FD1P3AX key_mem_14___i665 (.D(key_mem_0__127__N_6112[24]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [24])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i665.GSR = "ENABLED";
    FD1P3AX key_mem_14___i666 (.D(key_mem_0__127__N_6112[25]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [25])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i666.GSR = "ENABLED";
    FD1P3AX key_mem_14___i667 (.D(key_mem_0__127__N_6112[26]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [26])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i667.GSR = "ENABLED";
    FD1P3AX key_mem_14___i668 (.D(key_mem_0__127__N_6112[27]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [27])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i668.GSR = "ENABLED";
    FD1P3AX key_mem_14___i669 (.D(key_mem_0__127__N_6112[28]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [28])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i669.GSR = "ENABLED";
    FD1P3AX key_mem_14___i670 (.D(key_mem_0__127__N_6112[29]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [29])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i670.GSR = "ENABLED";
    FD1P3AX key_mem_14___i671 (.D(key_mem_0__127__N_6112[30]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [30])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i671.GSR = "ENABLED";
    FD1P3AX key_mem_14___i672 (.D(key_mem_0__127__N_6112[31]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [31])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i672.GSR = "ENABLED";
    FD1P3AX key_mem_14___i673 (.D(key_mem_0__127__N_6112[32]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [32])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i673.GSR = "ENABLED";
    FD1P3AX key_mem_14___i674 (.D(key_mem_0__127__N_6112[33]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [33])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i674.GSR = "ENABLED";
    FD1P3AX key_mem_14___i675 (.D(key_mem_0__127__N_6112[34]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [34])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i675.GSR = "ENABLED";
    FD1P3AX key_mem_14___i676 (.D(key_mem_0__127__N_6112[35]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [35])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i676.GSR = "ENABLED";
    FD1P3AX key_mem_14___i677 (.D(key_mem_0__127__N_6112[36]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [36])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i677.GSR = "ENABLED";
    FD1P3AX key_mem_14___i678 (.D(key_mem_0__127__N_6112[37]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [37])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i678.GSR = "ENABLED";
    FD1P3AX key_mem_14___i679 (.D(key_mem_0__127__N_6112[38]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [38])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i679.GSR = "ENABLED";
    FD1P3AX key_mem_14___i680 (.D(key_mem_0__127__N_6112[39]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [39])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i680.GSR = "ENABLED";
    FD1P3AX key_mem_14___i681 (.D(key_mem_0__127__N_6112[40]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [40])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i681.GSR = "ENABLED";
    FD1P3AX key_mem_14___i682 (.D(key_mem_0__127__N_6112[41]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [41])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i682.GSR = "ENABLED";
    FD1P3AX key_mem_14___i683 (.D(key_mem_0__127__N_6112[42]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [42])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i683.GSR = "ENABLED";
    FD1P3AX key_mem_14___i684 (.D(key_mem_0__127__N_6112[43]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [43])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i684.GSR = "ENABLED";
    FD1P3AX key_mem_14___i685 (.D(key_mem_0__127__N_6112[44]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [44])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i685.GSR = "ENABLED";
    FD1P3AX key_mem_14___i686 (.D(key_mem_0__127__N_6112[45]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [45])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i686.GSR = "ENABLED";
    FD1P3AX key_mem_14___i687 (.D(key_mem_0__127__N_6112[46]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [46])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i687.GSR = "ENABLED";
    FD1P3AX key_mem_14___i688 (.D(key_mem_0__127__N_6112[47]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [47])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i688.GSR = "ENABLED";
    FD1P3AX key_mem_14___i689 (.D(key_mem_0__127__N_6112[48]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [48])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i689.GSR = "ENABLED";
    FD1P3AX key_mem_14___i690 (.D(key_mem_0__127__N_6112[49]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [49])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i690.GSR = "ENABLED";
    FD1P3AX key_mem_14___i691 (.D(key_mem_0__127__N_6112[50]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [50])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i691.GSR = "ENABLED";
    FD1P3AX key_mem_14___i692 (.D(key_mem_0__127__N_6112[51]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [51])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i692.GSR = "ENABLED";
    FD1P3AX key_mem_14___i693 (.D(key_mem_0__127__N_6112[52]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [52])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i693.GSR = "ENABLED";
    FD1P3AX key_mem_14___i694 (.D(key_mem_0__127__N_6112[53]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [53])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i694.GSR = "ENABLED";
    FD1P3AX key_mem_14___i695 (.D(key_mem_0__127__N_6112[54]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [54])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i695.GSR = "ENABLED";
    FD1P3AX key_mem_14___i696 (.D(key_mem_0__127__N_6112[55]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [55])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i696.GSR = "ENABLED";
    FD1P3AX key_mem_14___i697 (.D(key_mem_0__127__N_6112[56]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [56])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i697.GSR = "ENABLED";
    FD1P3AX key_mem_14___i698 (.D(key_mem_0__127__N_6112[57]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [57])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i698.GSR = "ENABLED";
    FD1P3AX key_mem_14___i699 (.D(key_mem_0__127__N_6112[58]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [58])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i699.GSR = "ENABLED";
    FD1P3AX key_mem_14___i700 (.D(key_mem_0__127__N_6112[59]), .SP(clk_c_enable_1086), 
            .CK(clk_c), .Q(\key_mem[9] [59])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i700.GSR = "ENABLED";
    FD1P3AX key_mem_14___i701 (.D(key_mem_0__127__N_6112[60]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [60])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i701.GSR = "ENABLED";
    FD1P3AX key_mem_14___i702 (.D(key_mem_0__127__N_6112[61]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [61])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i702.GSR = "ENABLED";
    FD1P3AX key_mem_14___i703 (.D(key_mem_0__127__N_6112[62]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [62])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i703.GSR = "ENABLED";
    FD1P3AX key_mem_14___i704 (.D(key_mem_0__127__N_6112[63]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [63])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i704.GSR = "ENABLED";
    FD1P3AX key_mem_14___i705 (.D(key_mem_0__127__N_6112[64]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [64])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i705.GSR = "ENABLED";
    FD1P3AX key_mem_14___i706 (.D(key_mem_0__127__N_6112[65]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [65])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i706.GSR = "ENABLED";
    FD1P3AX key_mem_14___i707 (.D(key_mem_0__127__N_6112[66]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [66])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i707.GSR = "ENABLED";
    FD1P3AX key_mem_14___i708 (.D(key_mem_0__127__N_6112[67]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [67])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i708.GSR = "ENABLED";
    FD1P3AX key_mem_14___i709 (.D(key_mem_0__127__N_6112[68]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [68])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i709.GSR = "ENABLED";
    FD1P3AX key_mem_14___i710 (.D(key_mem_0__127__N_6112[69]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [69])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i710.GSR = "ENABLED";
    FD1P3AX key_mem_14___i711 (.D(key_mem_0__127__N_6112[70]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [70])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i711.GSR = "ENABLED";
    FD1P3AX key_mem_14___i712 (.D(key_mem_0__127__N_6112[71]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [71])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i712.GSR = "ENABLED";
    FD1P3AX key_mem_14___i713 (.D(key_mem_0__127__N_6112[72]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [72])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i713.GSR = "ENABLED";
    FD1P3AX key_mem_14___i714 (.D(key_mem_0__127__N_6112[73]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [73])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i714.GSR = "ENABLED";
    FD1P3AX key_mem_14___i715 (.D(key_mem_0__127__N_6112[74]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [74])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i715.GSR = "ENABLED";
    FD1P3AX key_mem_14___i716 (.D(key_mem_0__127__N_6112[75]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [75])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i716.GSR = "ENABLED";
    FD1P3AX key_mem_14___i717 (.D(key_mem_0__127__N_6112[76]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [76])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i717.GSR = "ENABLED";
    FD1P3AX key_mem_14___i718 (.D(key_mem_0__127__N_6112[77]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [77])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i718.GSR = "ENABLED";
    FD1P3AX key_mem_14___i719 (.D(key_mem_0__127__N_6112[78]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [78])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i719.GSR = "ENABLED";
    FD1P3AX key_mem_14___i720 (.D(key_mem_0__127__N_6112[79]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [79])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i720.GSR = "ENABLED";
    FD1P3AX key_mem_14___i721 (.D(key_mem_0__127__N_6112[80]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [80])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i721.GSR = "ENABLED";
    FD1P3AX key_mem_14___i722 (.D(key_mem_0__127__N_6112[81]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [81])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i722.GSR = "ENABLED";
    FD1P3AX key_mem_14___i723 (.D(key_mem_0__127__N_6112[82]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [82])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i723.GSR = "ENABLED";
    FD1P3AX key_mem_14___i724 (.D(key_mem_0__127__N_6112[83]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [83])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i724.GSR = "ENABLED";
    FD1P3AX key_mem_14___i725 (.D(key_mem_0__127__N_6112[84]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [84])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i725.GSR = "ENABLED";
    FD1P3AX key_mem_14___i726 (.D(key_mem_0__127__N_6112[85]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [85])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i726.GSR = "ENABLED";
    FD1P3AX key_mem_14___i727 (.D(key_mem_0__127__N_6112[86]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [86])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i727.GSR = "ENABLED";
    FD1P3AX key_mem_14___i728 (.D(key_mem_0__127__N_6112[87]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [87])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i728.GSR = "ENABLED";
    FD1P3AX key_mem_14___i729 (.D(key_mem_0__127__N_6112[88]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [88])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i729.GSR = "ENABLED";
    FD1P3AX key_mem_14___i730 (.D(key_mem_0__127__N_6112[89]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [89])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i730.GSR = "ENABLED";
    FD1P3AX key_mem_14___i731 (.D(key_mem_0__127__N_6112[90]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [90])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i731.GSR = "ENABLED";
    FD1P3AX key_mem_14___i732 (.D(key_mem_0__127__N_6112[91]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [91])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i732.GSR = "ENABLED";
    FD1P3AX key_mem_14___i733 (.D(key_mem_0__127__N_6112[92]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [92])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i733.GSR = "ENABLED";
    FD1P3AX key_mem_14___i734 (.D(key_mem_0__127__N_6112[93]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [93])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i734.GSR = "ENABLED";
    FD1P3AX key_mem_14___i735 (.D(key_mem_0__127__N_6112[94]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [94])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i735.GSR = "ENABLED";
    FD1P3AX key_mem_14___i736 (.D(key_mem_0__127__N_6112[95]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [95])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i736.GSR = "ENABLED";
    FD1P3AX key_mem_14___i737 (.D(key_mem_0__127__N_6112[96]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [96])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i737.GSR = "ENABLED";
    FD1P3AX key_mem_14___i738 (.D(key_mem_0__127__N_6112[97]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [97])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i738.GSR = "ENABLED";
    FD1P3AX key_mem_14___i739 (.D(key_mem_0__127__N_6112[98]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [98])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i739.GSR = "ENABLED";
    FD1P3AX key_mem_14___i740 (.D(key_mem_0__127__N_6112[99]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [99])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i740.GSR = "ENABLED";
    FD1P3AX key_mem_14___i741 (.D(key_mem_0__127__N_6112[100]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [100])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i741.GSR = "ENABLED";
    FD1P3AX key_mem_14___i742 (.D(key_mem_0__127__N_6112[101]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [101])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i742.GSR = "ENABLED";
    FD1P3AX key_mem_14___i743 (.D(key_mem_0__127__N_6112[102]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [102])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i743.GSR = "ENABLED";
    FD1P3AX key_mem_14___i744 (.D(key_mem_0__127__N_6112[103]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [103])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i744.GSR = "ENABLED";
    FD1P3AX key_mem_14___i745 (.D(key_mem_0__127__N_6112[104]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [104])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i745.GSR = "ENABLED";
    FD1P3AX key_mem_14___i746 (.D(key_mem_0__127__N_6112[105]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [105])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i746.GSR = "ENABLED";
    FD1P3AX key_mem_14___i747 (.D(key_mem_0__127__N_6112[106]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [106])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i747.GSR = "ENABLED";
    FD1P3AX key_mem_14___i748 (.D(key_mem_0__127__N_6112[107]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [107])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i748.GSR = "ENABLED";
    FD1P3AX key_mem_14___i749 (.D(key_mem_0__127__N_6112[108]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [108])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i749.GSR = "ENABLED";
    FD1P3AX key_mem_14___i750 (.D(key_mem_0__127__N_6112[109]), .SP(clk_c_enable_1136), 
            .CK(clk_c), .Q(\key_mem[9] [109])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i750.GSR = "ENABLED";
    FD1P3AX key_mem_14___i751 (.D(key_mem_0__127__N_6112[110]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[9] [110])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i751.GSR = "ENABLED";
    FD1P3AX key_mem_14___i752 (.D(key_mem_0__127__N_6112[111]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[9] [111])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i752.GSR = "ENABLED";
    FD1P3AX key_mem_14___i753 (.D(key_mem_0__127__N_6112[112]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[9] [112])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i753.GSR = "ENABLED";
    FD1P3AX key_mem_14___i754 (.D(key_mem_0__127__N_6112[113]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[9] [113])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i754.GSR = "ENABLED";
    FD1P3AX key_mem_14___i755 (.D(key_mem_0__127__N_6112[114]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[9] [114])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i755.GSR = "ENABLED";
    FD1P3AX key_mem_14___i756 (.D(key_mem_0__127__N_6112[115]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[9] [115])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i756.GSR = "ENABLED";
    FD1P3AX key_mem_14___i757 (.D(key_mem_0__127__N_6112[116]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[9] [116])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i757.GSR = "ENABLED";
    FD1P3AX key_mem_14___i758 (.D(key_mem_0__127__N_6112[117]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[9] [117])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i758.GSR = "ENABLED";
    FD1P3AX key_mem_14___i759 (.D(key_mem_0__127__N_6112[118]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[9] [118])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i759.GSR = "ENABLED";
    FD1P3AX key_mem_14___i760 (.D(key_mem_0__127__N_6112[119]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[9] [119])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i760.GSR = "ENABLED";
    FD1P3AX key_mem_14___i761 (.D(key_mem_0__127__N_6112[120]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[9] [120])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i761.GSR = "ENABLED";
    FD1P3AX key_mem_14___i762 (.D(key_mem_0__127__N_6112[121]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[9] [121])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i762.GSR = "ENABLED";
    FD1P3AX key_mem_14___i763 (.D(key_mem_0__127__N_6112[122]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[9] [122])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i763.GSR = "ENABLED";
    FD1P3AX key_mem_14___i764 (.D(key_mem_0__127__N_6112[123]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[9] [123])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i764.GSR = "ENABLED";
    FD1P3AX key_mem_14___i765 (.D(key_mem_0__127__N_6112[124]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[9] [124])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i765.GSR = "ENABLED";
    FD1P3AX key_mem_14___i766 (.D(key_mem_0__127__N_6112[125]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[9] [125])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i766.GSR = "ENABLED";
    FD1P3AX key_mem_14___i767 (.D(key_mem_0__127__N_6112[126]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[9] [126])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i767.GSR = "ENABLED";
    FD1P3AX key_mem_14___i768 (.D(key_mem_0__127__N_6112[127]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[9] [127])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i768.GSR = "ENABLED";
    FD1P3AX key_mem_14___i769 (.D(key_mem_0__127__N_5984[0]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[8] [0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i769.GSR = "ENABLED";
    FD1P3AX key_mem_14___i770 (.D(key_mem_0__127__N_5984[1]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[8] [1])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i770.GSR = "ENABLED";
    FD1P3AX key_mem_14___i771 (.D(key_mem_0__127__N_5984[2]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[8] [2])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i771.GSR = "ENABLED";
    FD1P3AX key_mem_14___i772 (.D(key_mem_0__127__N_5984[3]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[8] [3])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i772.GSR = "ENABLED";
    FD1P3AX key_mem_14___i773 (.D(key_mem_0__127__N_5984[4]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[8] [4])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i773.GSR = "ENABLED";
    FD1P3AX key_mem_14___i774 (.D(key_mem_0__127__N_5984[5]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[8] [5])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i774.GSR = "ENABLED";
    FD1P3AX key_mem_14___i775 (.D(key_mem_0__127__N_5984[6]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[8] [6])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i775.GSR = "ENABLED";
    FD1P3AX key_mem_14___i776 (.D(key_mem_0__127__N_5984[7]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[8] [7])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i776.GSR = "ENABLED";
    FD1P3AX key_mem_14___i777 (.D(key_mem_0__127__N_5984[8]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[8] [8])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i777.GSR = "ENABLED";
    FD1P3AX key_mem_14___i778 (.D(key_mem_0__127__N_5984[9]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[8] [9])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i778.GSR = "ENABLED";
    FD1P3AX key_mem_14___i779 (.D(key_mem_0__127__N_5984[10]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[8] [10])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i779.GSR = "ENABLED";
    FD1P3AX key_mem_14___i780 (.D(key_mem_0__127__N_5984[11]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[8] [11])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i780.GSR = "ENABLED";
    FD1P3AX key_mem_14___i781 (.D(key_mem_0__127__N_5984[12]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[8] [12])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i781.GSR = "ENABLED";
    FD1P3AX key_mem_14___i782 (.D(key_mem_0__127__N_5984[13]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[8] [13])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i782.GSR = "ENABLED";
    FD1P3AX key_mem_14___i783 (.D(key_mem_0__127__N_5984[14]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[8] [14])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i783.GSR = "ENABLED";
    FD1P3AX key_mem_14___i784 (.D(key_mem_0__127__N_5984[15]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[8] [15])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i784.GSR = "ENABLED";
    FD1P3AX key_mem_14___i785 (.D(key_mem_0__127__N_5984[16]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[8] [16])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i785.GSR = "ENABLED";
    FD1P3AX key_mem_14___i786 (.D(key_mem_0__127__N_5984[17]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[8] [17])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i786.GSR = "ENABLED";
    FD1P3AX key_mem_14___i787 (.D(key_mem_0__127__N_5984[18]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[8] [18])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i787.GSR = "ENABLED";
    FD1P3AX key_mem_14___i788 (.D(key_mem_0__127__N_5984[19]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[8] [19])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i788.GSR = "ENABLED";
    FD1P3AX key_mem_14___i789 (.D(key_mem_0__127__N_5984[20]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[8] [20])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i789.GSR = "ENABLED";
    FD1P3AX key_mem_14___i790 (.D(key_mem_0__127__N_5984[21]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[8] [21])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i790.GSR = "ENABLED";
    FD1P3AX key_mem_14___i791 (.D(key_mem_0__127__N_5984[22]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[8] [22])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i791.GSR = "ENABLED";
    FD1P3AX key_mem_14___i792 (.D(key_mem_0__127__N_5984[23]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[8] [23])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i792.GSR = "ENABLED";
    FD1P3AX key_mem_14___i793 (.D(key_mem_0__127__N_5984[24]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[8] [24])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i793.GSR = "ENABLED";
    FD1P3AX key_mem_14___i794 (.D(key_mem_0__127__N_5984[25]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[8] [25])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i794.GSR = "ENABLED";
    FD1P3AX key_mem_14___i795 (.D(key_mem_0__127__N_5984[26]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[8] [26])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i795.GSR = "ENABLED";
    FD1P3AX key_mem_14___i796 (.D(key_mem_0__127__N_5984[27]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[8] [27])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i796.GSR = "ENABLED";
    FD1P3AX key_mem_14___i797 (.D(key_mem_0__127__N_5984[28]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[8] [28])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i797.GSR = "ENABLED";
    FD1P3AX key_mem_14___i798 (.D(key_mem_0__127__N_5984[29]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[8] [29])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i798.GSR = "ENABLED";
    FD1P3AX key_mem_14___i799 (.D(key_mem_0__127__N_5984[30]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[8] [30])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i799.GSR = "ENABLED";
    FD1P3AX key_mem_14___i800 (.D(key_mem_0__127__N_5984[31]), .SP(clk_c_enable_1186), 
            .CK(clk_c), .Q(\key_mem[8] [31])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i800.GSR = "ENABLED";
    FD1P3AX key_mem_14___i801 (.D(key_mem_0__127__N_5984[32]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [32])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i801.GSR = "ENABLED";
    FD1P3AX key_mem_14___i802 (.D(key_mem_0__127__N_5984[33]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [33])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i802.GSR = "ENABLED";
    FD1P3AX key_mem_14___i803 (.D(key_mem_0__127__N_5984[34]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [34])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i803.GSR = "ENABLED";
    FD1P3AX key_mem_14___i804 (.D(key_mem_0__127__N_5984[35]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [35])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i804.GSR = "ENABLED";
    FD1P3AX key_mem_14___i805 (.D(key_mem_0__127__N_5984[36]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [36])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i805.GSR = "ENABLED";
    FD1P3AX key_mem_14___i806 (.D(key_mem_0__127__N_5984[37]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [37])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i806.GSR = "ENABLED";
    FD1P3AX key_mem_14___i807 (.D(key_mem_0__127__N_5984[38]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [38])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i807.GSR = "ENABLED";
    FD1P3AX key_mem_14___i808 (.D(key_mem_0__127__N_5984[39]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [39])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i808.GSR = "ENABLED";
    FD1P3AX key_mem_14___i809 (.D(key_mem_0__127__N_5984[40]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [40])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i809.GSR = "ENABLED";
    FD1P3AX key_mem_14___i810 (.D(key_mem_0__127__N_5984[41]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [41])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i810.GSR = "ENABLED";
    FD1P3AX key_mem_14___i811 (.D(key_mem_0__127__N_5984[42]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [42])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i811.GSR = "ENABLED";
    FD1P3AX key_mem_14___i812 (.D(key_mem_0__127__N_5984[43]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [43])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i812.GSR = "ENABLED";
    FD1P3AX key_mem_14___i813 (.D(key_mem_0__127__N_5984[44]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [44])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i813.GSR = "ENABLED";
    FD1P3AX key_mem_14___i814 (.D(key_mem_0__127__N_5984[45]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [45])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i814.GSR = "ENABLED";
    FD1P3AX key_mem_14___i815 (.D(key_mem_0__127__N_5984[46]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [46])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i815.GSR = "ENABLED";
    FD1P3AX key_mem_14___i816 (.D(key_mem_0__127__N_5984[47]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [47])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i816.GSR = "ENABLED";
    FD1P3AX key_mem_14___i817 (.D(key_mem_0__127__N_5984[48]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [48])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i817.GSR = "ENABLED";
    FD1P3AX key_mem_14___i818 (.D(key_mem_0__127__N_5984[49]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [49])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i818.GSR = "ENABLED";
    FD1P3AX key_mem_14___i819 (.D(key_mem_0__127__N_5984[50]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [50])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i819.GSR = "ENABLED";
    FD1P3AX key_mem_14___i820 (.D(key_mem_0__127__N_5984[51]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [51])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i820.GSR = "ENABLED";
    FD1P3AX key_mem_14___i821 (.D(key_mem_0__127__N_5984[52]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [52])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i821.GSR = "ENABLED";
    FD1P3AX key_mem_14___i822 (.D(key_mem_0__127__N_5984[53]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [53])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i822.GSR = "ENABLED";
    FD1P3AX key_mem_14___i823 (.D(key_mem_0__127__N_5984[54]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [54])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i823.GSR = "ENABLED";
    FD1P3AX key_mem_14___i824 (.D(key_mem_0__127__N_5984[55]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [55])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i824.GSR = "ENABLED";
    FD1P3AX key_mem_14___i825 (.D(key_mem_0__127__N_5984[56]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [56])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i825.GSR = "ENABLED";
    FD1P3AX key_mem_14___i826 (.D(key_mem_0__127__N_5984[57]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [57])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i826.GSR = "ENABLED";
    FD1P3AX key_mem_14___i827 (.D(key_mem_0__127__N_5984[58]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [58])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i827.GSR = "ENABLED";
    FD1P3AX key_mem_14___i828 (.D(key_mem_0__127__N_5984[59]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [59])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i828.GSR = "ENABLED";
    FD1P3AX key_mem_14___i829 (.D(key_mem_0__127__N_5984[60]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [60])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i829.GSR = "ENABLED";
    FD1P3AX key_mem_14___i830 (.D(key_mem_0__127__N_5984[61]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [61])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i830.GSR = "ENABLED";
    FD1P3AX key_mem_14___i831 (.D(key_mem_0__127__N_5984[62]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [62])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i831.GSR = "ENABLED";
    FD1P3AX key_mem_14___i832 (.D(key_mem_0__127__N_5984[63]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [63])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i832.GSR = "ENABLED";
    FD1P3AX key_mem_14___i833 (.D(key_mem_0__127__N_5984[64]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [64])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i833.GSR = "ENABLED";
    FD1P3AX key_mem_14___i834 (.D(key_mem_0__127__N_5984[65]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [65])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i834.GSR = "ENABLED";
    FD1P3AX key_mem_14___i835 (.D(key_mem_0__127__N_5984[66]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [66])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i835.GSR = "ENABLED";
    FD1P3AX key_mem_14___i836 (.D(key_mem_0__127__N_5984[67]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [67])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i836.GSR = "ENABLED";
    FD1P3AX key_mem_14___i837 (.D(key_mem_0__127__N_5984[68]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [68])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i837.GSR = "ENABLED";
    FD1P3AX key_mem_14___i838 (.D(key_mem_0__127__N_5984[69]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [69])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i838.GSR = "ENABLED";
    FD1P3AX key_mem_14___i839 (.D(key_mem_0__127__N_5984[70]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [70])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i839.GSR = "ENABLED";
    FD1P3AX key_mem_14___i840 (.D(key_mem_0__127__N_5984[71]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [71])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i840.GSR = "ENABLED";
    FD1P3AX key_mem_14___i841 (.D(key_mem_0__127__N_5984[72]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [72])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i841.GSR = "ENABLED";
    FD1P3AX key_mem_14___i842 (.D(key_mem_0__127__N_5984[73]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [73])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i842.GSR = "ENABLED";
    FD1P3AX key_mem_14___i843 (.D(key_mem_0__127__N_5984[74]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [74])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i843.GSR = "ENABLED";
    FD1P3AX key_mem_14___i844 (.D(key_mem_0__127__N_5984[75]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [75])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i844.GSR = "ENABLED";
    FD1P3AX key_mem_14___i845 (.D(key_mem_0__127__N_5984[76]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [76])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i845.GSR = "ENABLED";
    FD1P3AX key_mem_14___i846 (.D(key_mem_0__127__N_5984[77]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [77])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i846.GSR = "ENABLED";
    FD1P3AX key_mem_14___i847 (.D(key_mem_0__127__N_5984[78]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [78])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i847.GSR = "ENABLED";
    FD1P3AX key_mem_14___i848 (.D(key_mem_0__127__N_5984[79]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [79])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i848.GSR = "ENABLED";
    FD1P3AX key_mem_14___i849 (.D(key_mem_0__127__N_5984[80]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [80])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i849.GSR = "ENABLED";
    FD1P3AX key_mem_14___i850 (.D(key_mem_0__127__N_5984[81]), .SP(clk_c_enable_1236), 
            .CK(clk_c), .Q(\key_mem[8] [81])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i850.GSR = "ENABLED";
    FD1P3AX key_mem_14___i851 (.D(key_mem_0__127__N_5984[82]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[8] [82])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i851.GSR = "ENABLED";
    FD1P3AX key_mem_14___i852 (.D(key_mem_0__127__N_5984[83]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[8] [83])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i852.GSR = "ENABLED";
    FD1P3AX key_mem_14___i853 (.D(key_mem_0__127__N_5984[84]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[8] [84])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i853.GSR = "ENABLED";
    FD1P3AX key_mem_14___i854 (.D(key_mem_0__127__N_5984[85]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[8] [85])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i854.GSR = "ENABLED";
    FD1P3AX key_mem_14___i855 (.D(key_mem_0__127__N_5984[86]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[8] [86])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i855.GSR = "ENABLED";
    FD1P3AX key_mem_14___i856 (.D(key_mem_0__127__N_5984[87]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[8] [87])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i856.GSR = "ENABLED";
    FD1P3AX key_mem_14___i857 (.D(key_mem_0__127__N_5984[88]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[8] [88])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i857.GSR = "ENABLED";
    FD1P3AX key_mem_14___i858 (.D(key_mem_0__127__N_5984[89]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[8] [89])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i858.GSR = "ENABLED";
    FD1P3AX key_mem_14___i859 (.D(key_mem_0__127__N_5984[90]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[8] [90])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i859.GSR = "ENABLED";
    FD1P3AX key_mem_14___i860 (.D(key_mem_0__127__N_5984[91]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[8] [91])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i860.GSR = "ENABLED";
    FD1P3AX key_mem_14___i861 (.D(key_mem_0__127__N_5984[92]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[8] [92])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i861.GSR = "ENABLED";
    FD1P3AX key_mem_14___i862 (.D(key_mem_0__127__N_5984[93]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[8] [93])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i862.GSR = "ENABLED";
    FD1P3AX key_mem_14___i863 (.D(key_mem_0__127__N_5984[94]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[8] [94])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i863.GSR = "ENABLED";
    FD1P3AX key_mem_14___i864 (.D(key_mem_0__127__N_5984[95]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[8] [95])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i864.GSR = "ENABLED";
    FD1P3AX key_mem_14___i865 (.D(key_mem_0__127__N_5984[96]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[8] [96])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i865.GSR = "ENABLED";
    FD1P3AX key_mem_14___i866 (.D(key_mem_0__127__N_5984[97]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[8] [97])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i866.GSR = "ENABLED";
    FD1P3AX key_mem_14___i867 (.D(key_mem_0__127__N_5984[98]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[8] [98])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i867.GSR = "ENABLED";
    FD1P3AX key_mem_14___i868 (.D(key_mem_0__127__N_5984[99]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[8] [99])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i868.GSR = "ENABLED";
    FD1P3AX key_mem_14___i869 (.D(key_mem_0__127__N_5984[100]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[8] [100])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i869.GSR = "ENABLED";
    FD1P3AX key_mem_14___i870 (.D(key_mem_0__127__N_5984[101]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[8] [101])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i870.GSR = "ENABLED";
    FD1P3AX key_mem_14___i871 (.D(key_mem_0__127__N_5984[102]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[8] [102])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i871.GSR = "ENABLED";
    FD1P3AX key_mem_14___i872 (.D(key_mem_0__127__N_5984[103]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[8] [103])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i872.GSR = "ENABLED";
    FD1P3AX key_mem_14___i873 (.D(key_mem_0__127__N_5984[104]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[8] [104])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i873.GSR = "ENABLED";
    FD1P3AX key_mem_14___i874 (.D(key_mem_0__127__N_5984[105]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[8] [105])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i874.GSR = "ENABLED";
    FD1P3AX key_mem_14___i875 (.D(key_mem_0__127__N_5984[106]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[8] [106])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i875.GSR = "ENABLED";
    FD1P3AX key_mem_14___i876 (.D(key_mem_0__127__N_5984[107]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[8] [107])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i876.GSR = "ENABLED";
    FD1P3AX key_mem_14___i877 (.D(key_mem_0__127__N_5984[108]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[8] [108])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i877.GSR = "ENABLED";
    FD1P3AX key_mem_14___i878 (.D(key_mem_0__127__N_5984[109]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[8] [109])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i878.GSR = "ENABLED";
    FD1P3AX key_mem_14___i879 (.D(key_mem_0__127__N_5984[110]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[8] [110])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i879.GSR = "ENABLED";
    FD1P3AX key_mem_14___i880 (.D(key_mem_0__127__N_5984[111]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[8] [111])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i880.GSR = "ENABLED";
    FD1P3AX key_mem_14___i881 (.D(key_mem_0__127__N_5984[112]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[8] [112])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i881.GSR = "ENABLED";
    FD1P3AX key_mem_14___i882 (.D(key_mem_0__127__N_5984[113]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[8] [113])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i882.GSR = "ENABLED";
    FD1P3AX key_mem_14___i883 (.D(key_mem_0__127__N_5984[114]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[8] [114])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i883.GSR = "ENABLED";
    FD1P3AX key_mem_14___i884 (.D(key_mem_0__127__N_5984[115]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[8] [115])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i884.GSR = "ENABLED";
    FD1P3AX key_mem_14___i885 (.D(key_mem_0__127__N_5984[116]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[8] [116])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i885.GSR = "ENABLED";
    FD1P3AX key_mem_14___i886 (.D(key_mem_0__127__N_5984[117]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[8] [117])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i886.GSR = "ENABLED";
    FD1P3AX key_mem_14___i887 (.D(key_mem_0__127__N_5984[118]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[8] [118])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i887.GSR = "ENABLED";
    FD1P3AX key_mem_14___i888 (.D(key_mem_0__127__N_5984[119]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[8] [119])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i888.GSR = "ENABLED";
    FD1P3AX key_mem_14___i889 (.D(key_mem_0__127__N_5984[120]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[8] [120])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i889.GSR = "ENABLED";
    FD1P3AX key_mem_14___i890 (.D(key_mem_0__127__N_5984[121]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[8] [121])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i890.GSR = "ENABLED";
    FD1P3AX key_mem_14___i891 (.D(key_mem_0__127__N_5984[122]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[8] [122])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i891.GSR = "ENABLED";
    FD1P3AX key_mem_14___i892 (.D(key_mem_0__127__N_5984[123]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[8] [123])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i892.GSR = "ENABLED";
    FD1P3AX key_mem_14___i893 (.D(key_mem_0__127__N_5984[124]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[8] [124])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i893.GSR = "ENABLED";
    FD1P3AX key_mem_14___i894 (.D(key_mem_0__127__N_5984[125]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[8] [125])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i894.GSR = "ENABLED";
    FD1P3AX key_mem_14___i895 (.D(key_mem_0__127__N_5984[126]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[8] [126])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i895.GSR = "ENABLED";
    FD1P3AX key_mem_14___i896 (.D(key_mem_0__127__N_5984[127]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[8] [127])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i896.GSR = "ENABLED";
    FD1P3AX key_mem_14___i897 (.D(key_mem_0__127__N_5856[0]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[7] [0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i897.GSR = "ENABLED";
    FD1P3AX key_mem_14___i898 (.D(key_mem_0__127__N_5856[1]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[7] [1])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i898.GSR = "ENABLED";
    FD1P3AX key_mem_14___i899 (.D(key_mem_0__127__N_5856[2]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[7] [2])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i899.GSR = "ENABLED";
    FD1P3AX key_mem_14___i900 (.D(key_mem_0__127__N_5856[3]), .SP(clk_c_enable_1286), 
            .CK(clk_c), .Q(\key_mem[7] [3])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i900.GSR = "ENABLED";
    FD1P3AX key_mem_14___i901 (.D(key_mem_0__127__N_5856[4]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [4])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i901.GSR = "ENABLED";
    FD1P3AX key_mem_14___i902 (.D(key_mem_0__127__N_5856[5]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [5])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i902.GSR = "ENABLED";
    FD1P3AX key_mem_14___i903 (.D(key_mem_0__127__N_5856[6]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [6])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i903.GSR = "ENABLED";
    FD1P3AX key_mem_14___i904 (.D(key_mem_0__127__N_5856[7]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [7])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i904.GSR = "ENABLED";
    FD1P3AX key_mem_14___i905 (.D(key_mem_0__127__N_5856[8]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [8])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i905.GSR = "ENABLED";
    FD1P3AX key_mem_14___i906 (.D(key_mem_0__127__N_5856[9]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [9])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i906.GSR = "ENABLED";
    FD1P3AX key_mem_14___i907 (.D(key_mem_0__127__N_5856[10]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [10])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i907.GSR = "ENABLED";
    FD1P3AX key_mem_14___i908 (.D(key_mem_0__127__N_5856[11]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [11])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i908.GSR = "ENABLED";
    FD1P3AX key_mem_14___i909 (.D(key_mem_0__127__N_5856[12]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [12])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i909.GSR = "ENABLED";
    FD1P3AX key_mem_14___i910 (.D(key_mem_0__127__N_5856[13]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [13])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i910.GSR = "ENABLED";
    FD1P3AX key_mem_14___i911 (.D(key_mem_0__127__N_5856[14]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [14])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i911.GSR = "ENABLED";
    FD1P3AX key_mem_14___i912 (.D(key_mem_0__127__N_5856[15]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [15])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i912.GSR = "ENABLED";
    FD1P3AX key_mem_14___i913 (.D(key_mem_0__127__N_5856[16]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [16])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i913.GSR = "ENABLED";
    FD1P3AX key_mem_14___i914 (.D(key_mem_0__127__N_5856[17]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [17])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i914.GSR = "ENABLED";
    FD1P3AX key_mem_14___i915 (.D(key_mem_0__127__N_5856[18]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [18])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i915.GSR = "ENABLED";
    FD1P3AX key_mem_14___i916 (.D(key_mem_0__127__N_5856[19]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [19])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i916.GSR = "ENABLED";
    FD1P3AX key_mem_14___i917 (.D(key_mem_0__127__N_5856[20]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [20])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i917.GSR = "ENABLED";
    FD1P3AX key_mem_14___i918 (.D(key_mem_0__127__N_5856[21]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [21])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i918.GSR = "ENABLED";
    FD1P3AX key_mem_14___i919 (.D(key_mem_0__127__N_5856[22]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [22])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i919.GSR = "ENABLED";
    FD1P3AX key_mem_14___i920 (.D(key_mem_0__127__N_5856[23]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [23])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i920.GSR = "ENABLED";
    FD1P3AX key_mem_14___i921 (.D(key_mem_0__127__N_5856[24]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [24])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i921.GSR = "ENABLED";
    FD1P3AX key_mem_14___i922 (.D(key_mem_0__127__N_5856[25]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [25])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i922.GSR = "ENABLED";
    FD1P3AX key_mem_14___i923 (.D(key_mem_0__127__N_5856[26]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [26])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i923.GSR = "ENABLED";
    FD1P3AX key_mem_14___i924 (.D(key_mem_0__127__N_5856[27]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [27])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i924.GSR = "ENABLED";
    FD1P3AX key_mem_14___i925 (.D(key_mem_0__127__N_5856[28]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [28])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i925.GSR = "ENABLED";
    FD1P3AX key_mem_14___i926 (.D(key_mem_0__127__N_5856[29]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [29])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i926.GSR = "ENABLED";
    FD1P3AX key_mem_14___i927 (.D(key_mem_0__127__N_5856[30]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [30])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i927.GSR = "ENABLED";
    FD1P3AX key_mem_14___i928 (.D(key_mem_0__127__N_5856[31]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [31])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i928.GSR = "ENABLED";
    FD1P3AX key_mem_14___i929 (.D(key_mem_0__127__N_5856[32]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [32])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i929.GSR = "ENABLED";
    FD1P3AX key_mem_14___i930 (.D(key_mem_0__127__N_5856[33]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [33])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i930.GSR = "ENABLED";
    FD1P3AX key_mem_14___i931 (.D(key_mem_0__127__N_5856[34]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [34])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i931.GSR = "ENABLED";
    FD1P3AX key_mem_14___i932 (.D(key_mem_0__127__N_5856[35]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [35])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i932.GSR = "ENABLED";
    FD1P3AX key_mem_14___i933 (.D(key_mem_0__127__N_5856[36]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [36])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i933.GSR = "ENABLED";
    FD1P3AX key_mem_14___i934 (.D(key_mem_0__127__N_5856[37]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [37])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i934.GSR = "ENABLED";
    FD1P3AX key_mem_14___i935 (.D(key_mem_0__127__N_5856[38]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [38])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i935.GSR = "ENABLED";
    FD1P3AX key_mem_14___i936 (.D(key_mem_0__127__N_5856[39]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [39])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i936.GSR = "ENABLED";
    FD1P3AX key_mem_14___i937 (.D(key_mem_0__127__N_5856[40]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [40])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i937.GSR = "ENABLED";
    FD1P3AX key_mem_14___i938 (.D(key_mem_0__127__N_5856[41]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [41])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i938.GSR = "ENABLED";
    FD1P3AX key_mem_14___i939 (.D(key_mem_0__127__N_5856[42]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [42])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i939.GSR = "ENABLED";
    FD1P3AX key_mem_14___i940 (.D(key_mem_0__127__N_5856[43]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [43])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i940.GSR = "ENABLED";
    FD1P3AX key_mem_14___i941 (.D(key_mem_0__127__N_5856[44]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [44])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i941.GSR = "ENABLED";
    FD1P3AX key_mem_14___i942 (.D(key_mem_0__127__N_5856[45]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [45])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i942.GSR = "ENABLED";
    FD1P3AX key_mem_14___i943 (.D(key_mem_0__127__N_5856[46]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [46])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i943.GSR = "ENABLED";
    FD1P3AX key_mem_14___i944 (.D(key_mem_0__127__N_5856[47]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [47])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i944.GSR = "ENABLED";
    FD1P3AX key_mem_14___i945 (.D(key_mem_0__127__N_5856[48]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [48])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i945.GSR = "ENABLED";
    FD1P3AX key_mem_14___i946 (.D(key_mem_0__127__N_5856[49]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [49])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i946.GSR = "ENABLED";
    FD1P3AX key_mem_14___i947 (.D(key_mem_0__127__N_5856[50]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [50])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i947.GSR = "ENABLED";
    FD1P3AX key_mem_14___i948 (.D(key_mem_0__127__N_5856[51]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [51])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i948.GSR = "ENABLED";
    FD1P3AX key_mem_14___i949 (.D(key_mem_0__127__N_5856[52]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [52])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i949.GSR = "ENABLED";
    FD1P3AX key_mem_14___i950 (.D(key_mem_0__127__N_5856[53]), .SP(clk_c_enable_1336), 
            .CK(clk_c), .Q(\key_mem[7] [53])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i950.GSR = "ENABLED";
    FD1P3AX key_mem_14___i951 (.D(key_mem_0__127__N_5856[54]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [54])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i951.GSR = "ENABLED";
    FD1P3AX key_mem_14___i952 (.D(key_mem_0__127__N_5856[55]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [55])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i952.GSR = "ENABLED";
    FD1P3AX key_mem_14___i953 (.D(key_mem_0__127__N_5856[56]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [56])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i953.GSR = "ENABLED";
    FD1P3AX key_mem_14___i954 (.D(key_mem_0__127__N_5856[57]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [57])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i954.GSR = "ENABLED";
    FD1P3AX key_mem_14___i955 (.D(key_mem_0__127__N_5856[58]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [58])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i955.GSR = "ENABLED";
    FD1P3AX key_mem_14___i956 (.D(key_mem_0__127__N_5856[59]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [59])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i956.GSR = "ENABLED";
    FD1P3AX key_mem_14___i957 (.D(key_mem_0__127__N_5856[60]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [60])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i957.GSR = "ENABLED";
    FD1P3AX key_mem_14___i958 (.D(key_mem_0__127__N_5856[61]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [61])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i958.GSR = "ENABLED";
    FD1P3AX key_mem_14___i959 (.D(key_mem_0__127__N_5856[62]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [62])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i959.GSR = "ENABLED";
    FD1P3AX key_mem_14___i960 (.D(key_mem_0__127__N_5856[63]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [63])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i960.GSR = "ENABLED";
    FD1P3AX key_mem_14___i961 (.D(key_mem_0__127__N_5856[64]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [64])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i961.GSR = "ENABLED";
    FD1P3AX key_mem_14___i962 (.D(key_mem_0__127__N_5856[65]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [65])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i962.GSR = "ENABLED";
    FD1P3AX key_mem_14___i963 (.D(key_mem_0__127__N_5856[66]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [66])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i963.GSR = "ENABLED";
    FD1P3AX key_mem_14___i964 (.D(key_mem_0__127__N_5856[67]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [67])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i964.GSR = "ENABLED";
    FD1P3AX key_mem_14___i965 (.D(key_mem_0__127__N_5856[68]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [68])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i965.GSR = "ENABLED";
    FD1P3AX key_mem_14___i966 (.D(key_mem_0__127__N_5856[69]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [69])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i966.GSR = "ENABLED";
    FD1P3AX key_mem_14___i967 (.D(key_mem_0__127__N_5856[70]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [70])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i967.GSR = "ENABLED";
    FD1P3AX key_mem_14___i968 (.D(key_mem_0__127__N_5856[71]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [71])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i968.GSR = "ENABLED";
    FD1P3AX key_mem_14___i969 (.D(key_mem_0__127__N_5856[72]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [72])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i969.GSR = "ENABLED";
    FD1P3AX key_mem_14___i970 (.D(key_mem_0__127__N_5856[73]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [73])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i970.GSR = "ENABLED";
    FD1P3AX key_mem_14___i971 (.D(key_mem_0__127__N_5856[74]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [74])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i971.GSR = "ENABLED";
    FD1P3AX key_mem_14___i972 (.D(key_mem_0__127__N_5856[75]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [75])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i972.GSR = "ENABLED";
    FD1P3AX key_mem_14___i973 (.D(key_mem_0__127__N_5856[76]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [76])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i973.GSR = "ENABLED";
    FD1P3AX key_mem_14___i974 (.D(key_mem_0__127__N_5856[77]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [77])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i974.GSR = "ENABLED";
    FD1P3AX key_mem_14___i975 (.D(key_mem_0__127__N_5856[78]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [78])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i975.GSR = "ENABLED";
    FD1P3AX key_mem_14___i976 (.D(key_mem_0__127__N_5856[79]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [79])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i976.GSR = "ENABLED";
    FD1P3AX key_mem_14___i977 (.D(key_mem_0__127__N_5856[80]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [80])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i977.GSR = "ENABLED";
    FD1P3AX key_mem_14___i978 (.D(key_mem_0__127__N_5856[81]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [81])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i978.GSR = "ENABLED";
    FD1P3AX key_mem_14___i979 (.D(key_mem_0__127__N_5856[82]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [82])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i979.GSR = "ENABLED";
    FD1P3AX key_mem_14___i980 (.D(key_mem_0__127__N_5856[83]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [83])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i980.GSR = "ENABLED";
    FD1P3AX key_mem_14___i981 (.D(key_mem_0__127__N_5856[84]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [84])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i981.GSR = "ENABLED";
    FD1P3AX key_mem_14___i982 (.D(key_mem_0__127__N_5856[85]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [85])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i982.GSR = "ENABLED";
    FD1P3AX key_mem_14___i983 (.D(key_mem_0__127__N_5856[86]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [86])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i983.GSR = "ENABLED";
    FD1P3AX key_mem_14___i984 (.D(key_mem_0__127__N_5856[87]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [87])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i984.GSR = "ENABLED";
    FD1P3AX key_mem_14___i985 (.D(key_mem_0__127__N_5856[88]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [88])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i985.GSR = "ENABLED";
    FD1P3AX key_mem_14___i986 (.D(key_mem_0__127__N_5856[89]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [89])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i986.GSR = "ENABLED";
    FD1P3AX key_mem_14___i987 (.D(key_mem_0__127__N_5856[90]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [90])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i987.GSR = "ENABLED";
    FD1P3AX key_mem_14___i988 (.D(key_mem_0__127__N_5856[91]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [91])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i988.GSR = "ENABLED";
    FD1P3AX key_mem_14___i989 (.D(key_mem_0__127__N_5856[92]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [92])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i989.GSR = "ENABLED";
    FD1P3AX key_mem_14___i990 (.D(key_mem_0__127__N_5856[93]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [93])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i990.GSR = "ENABLED";
    FD1P3AX key_mem_14___i991 (.D(key_mem_0__127__N_5856[94]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [94])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i991.GSR = "ENABLED";
    FD1P3AX key_mem_14___i992 (.D(key_mem_0__127__N_5856[95]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [95])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i992.GSR = "ENABLED";
    FD1P3AX key_mem_14___i993 (.D(key_mem_0__127__N_5856[96]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [96])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i993.GSR = "ENABLED";
    FD1P3AX key_mem_14___i994 (.D(key_mem_0__127__N_5856[97]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [97])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i994.GSR = "ENABLED";
    FD1P3AX key_mem_14___i995 (.D(key_mem_0__127__N_5856[98]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [98])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i995.GSR = "ENABLED";
    FD1P3AX key_mem_14___i996 (.D(key_mem_0__127__N_5856[99]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [99])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i996.GSR = "ENABLED";
    FD1P3AX key_mem_14___i997 (.D(key_mem_0__127__N_5856[100]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [100])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i997.GSR = "ENABLED";
    FD1P3AX key_mem_14___i998 (.D(key_mem_0__127__N_5856[101]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [101])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i998.GSR = "ENABLED";
    FD1P3AX key_mem_14___i999 (.D(key_mem_0__127__N_5856[102]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [102])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i999.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1000 (.D(key_mem_0__127__N_5856[103]), .SP(clk_c_enable_1386), 
            .CK(clk_c), .Q(\key_mem[7] [103])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1000.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1001 (.D(key_mem_0__127__N_5856[104]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[7] [104])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1001.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1002 (.D(key_mem_0__127__N_5856[105]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[7] [105])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1002.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1003 (.D(key_mem_0__127__N_5856[106]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[7] [106])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1003.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1004 (.D(key_mem_0__127__N_5856[107]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[7] [107])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1004.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1005 (.D(key_mem_0__127__N_5856[108]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[7] [108])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1005.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1006 (.D(key_mem_0__127__N_5856[109]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[7] [109])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1006.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1007 (.D(key_mem_0__127__N_5856[110]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[7] [110])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1007.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1008 (.D(key_mem_0__127__N_5856[111]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[7] [111])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1008.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1009 (.D(key_mem_0__127__N_5856[112]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[7] [112])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1009.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1010 (.D(key_mem_0__127__N_5856[113]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[7] [113])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1010.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1011 (.D(key_mem_0__127__N_5856[114]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[7] [114])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1011.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1012 (.D(key_mem_0__127__N_5856[115]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[7] [115])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1012.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1013 (.D(key_mem_0__127__N_5856[116]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[7] [116])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1013.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1014 (.D(key_mem_0__127__N_5856[117]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[7] [117])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1014.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1015 (.D(key_mem_0__127__N_5856[118]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[7] [118])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1015.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1016 (.D(key_mem_0__127__N_5856[119]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[7] [119])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1016.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1017 (.D(key_mem_0__127__N_5856[120]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[7] [120])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1017.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1018 (.D(key_mem_0__127__N_5856[121]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[7] [121])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1018.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1019 (.D(key_mem_0__127__N_5856[122]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[7] [122])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1019.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1020 (.D(key_mem_0__127__N_5856[123]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[7] [123])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1020.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1021 (.D(key_mem_0__127__N_5856[124]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[7] [124])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1021.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1022 (.D(key_mem_0__127__N_5856[125]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[7] [125])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1022.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1023 (.D(key_mem_0__127__N_5856[126]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[7] [126])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1023.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1024 (.D(key_mem_0__127__N_5856[127]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[7] [127])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1024.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1025 (.D(key_mem_0__127__N_5728[0]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[6] [0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1025.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1026 (.D(key_mem_0__127__N_5728[1]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[6] [1])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1026.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1027 (.D(key_mem_0__127__N_5728[2]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[6] [2])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1027.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1028 (.D(key_mem_0__127__N_5728[3]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[6] [3])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1028.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1029 (.D(key_mem_0__127__N_5728[4]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[6] [4])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1029.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1030 (.D(key_mem_0__127__N_5728[5]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[6] [5])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1030.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1031 (.D(key_mem_0__127__N_5728[6]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[6] [6])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1031.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1032 (.D(key_mem_0__127__N_5728[7]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[6] [7])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1032.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1033 (.D(key_mem_0__127__N_5728[8]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[6] [8])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1033.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1034 (.D(key_mem_0__127__N_5728[9]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[6] [9])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1034.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1035 (.D(key_mem_0__127__N_5728[10]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[6] [10])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1035.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1036 (.D(key_mem_0__127__N_5728[11]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[6] [11])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1036.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1037 (.D(key_mem_0__127__N_5728[12]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[6] [12])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1037.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1038 (.D(key_mem_0__127__N_5728[13]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[6] [13])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1038.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1039 (.D(key_mem_0__127__N_5728[14]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[6] [14])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1039.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1040 (.D(key_mem_0__127__N_5728[15]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[6] [15])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1040.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1041 (.D(key_mem_0__127__N_5728[16]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[6] [16])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1041.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1042 (.D(key_mem_0__127__N_5728[17]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[6] [17])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1042.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1043 (.D(key_mem_0__127__N_5728[18]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[6] [18])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1043.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1044 (.D(key_mem_0__127__N_5728[19]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[6] [19])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1044.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1045 (.D(key_mem_0__127__N_5728[20]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[6] [20])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1045.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1046 (.D(key_mem_0__127__N_5728[21]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[6] [21])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1046.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1047 (.D(key_mem_0__127__N_5728[22]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[6] [22])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1047.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1048 (.D(key_mem_0__127__N_5728[23]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[6] [23])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1048.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1049 (.D(key_mem_0__127__N_5728[24]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[6] [24])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1049.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1050 (.D(key_mem_0__127__N_5728[25]), .SP(clk_c_enable_1436), 
            .CK(clk_c), .Q(\key_mem[6] [25])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1050.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1051 (.D(key_mem_0__127__N_5728[26]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [26])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1051.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1052 (.D(key_mem_0__127__N_5728[27]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [27])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1052.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1053 (.D(key_mem_0__127__N_5728[28]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [28])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1053.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1054 (.D(key_mem_0__127__N_5728[29]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [29])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1054.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1055 (.D(key_mem_0__127__N_5728[30]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [30])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1055.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1056 (.D(key_mem_0__127__N_5728[31]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [31])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1056.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1057 (.D(key_mem_0__127__N_5728[32]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [32])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1057.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1058 (.D(key_mem_0__127__N_5728[33]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [33])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1058.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1059 (.D(key_mem_0__127__N_5728[34]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [34])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1059.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1060 (.D(key_mem_0__127__N_5728[35]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [35])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1060.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1061 (.D(key_mem_0__127__N_5728[36]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [36])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1061.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1062 (.D(key_mem_0__127__N_5728[37]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [37])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1062.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1063 (.D(key_mem_0__127__N_5728[38]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [38])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1063.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1064 (.D(key_mem_0__127__N_5728[39]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [39])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1064.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1065 (.D(key_mem_0__127__N_5728[40]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [40])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1065.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1066 (.D(key_mem_0__127__N_5728[41]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [41])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1066.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1067 (.D(key_mem_0__127__N_5728[42]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [42])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1067.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1068 (.D(key_mem_0__127__N_5728[43]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [43])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1068.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1069 (.D(key_mem_0__127__N_5728[44]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [44])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1069.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1070 (.D(key_mem_0__127__N_5728[45]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [45])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1070.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1071 (.D(key_mem_0__127__N_5728[46]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [46])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1071.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1072 (.D(key_mem_0__127__N_5728[47]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [47])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1072.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1073 (.D(key_mem_0__127__N_5728[48]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [48])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1073.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1074 (.D(key_mem_0__127__N_5728[49]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [49])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1074.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1075 (.D(key_mem_0__127__N_5728[50]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [50])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1075.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1076 (.D(key_mem_0__127__N_5728[51]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [51])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1076.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1077 (.D(key_mem_0__127__N_5728[52]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [52])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1077.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1078 (.D(key_mem_0__127__N_5728[53]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [53])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1078.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1079 (.D(key_mem_0__127__N_5728[54]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [54])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1079.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1080 (.D(key_mem_0__127__N_5728[55]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [55])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1080.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1081 (.D(key_mem_0__127__N_5728[56]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [56])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1081.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1082 (.D(key_mem_0__127__N_5728[57]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [57])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1082.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1083 (.D(key_mem_0__127__N_5728[58]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [58])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1083.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1084 (.D(key_mem_0__127__N_5728[59]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [59])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1084.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1085 (.D(key_mem_0__127__N_5728[60]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [60])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1085.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1086 (.D(key_mem_0__127__N_5728[61]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [61])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1086.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1087 (.D(key_mem_0__127__N_5728[62]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [62])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1087.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1088 (.D(key_mem_0__127__N_5728[63]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [63])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1088.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1089 (.D(key_mem_0__127__N_5728[64]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [64])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1089.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1090 (.D(key_mem_0__127__N_5728[65]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [65])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1090.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1091 (.D(key_mem_0__127__N_5728[66]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [66])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1091.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1092 (.D(key_mem_0__127__N_5728[67]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [67])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1092.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1093 (.D(key_mem_0__127__N_5728[68]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [68])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1093.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1094 (.D(key_mem_0__127__N_5728[69]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [69])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1094.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1095 (.D(key_mem_0__127__N_5728[70]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [70])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1095.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1096 (.D(key_mem_0__127__N_5728[71]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [71])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1096.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1097 (.D(key_mem_0__127__N_5728[72]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [72])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1097.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1098 (.D(key_mem_0__127__N_5728[73]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [73])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1098.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1099 (.D(key_mem_0__127__N_5728[74]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [74])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1099.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1100 (.D(key_mem_0__127__N_5728[75]), .SP(clk_c_enable_1486), 
            .CK(clk_c), .Q(\key_mem[6] [75])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1100.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1101 (.D(key_mem_0__127__N_5728[76]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [76])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1101.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1102 (.D(key_mem_0__127__N_5728[77]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [77])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1102.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1103 (.D(key_mem_0__127__N_5728[78]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [78])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1103.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1104 (.D(key_mem_0__127__N_5728[79]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [79])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1104.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1105 (.D(key_mem_0__127__N_5728[80]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [80])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1105.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1106 (.D(key_mem_0__127__N_5728[81]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [81])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1106.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1107 (.D(key_mem_0__127__N_5728[82]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [82])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1107.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1108 (.D(key_mem_0__127__N_5728[83]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [83])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1108.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1109 (.D(key_mem_0__127__N_5728[84]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [84])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1109.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1110 (.D(key_mem_0__127__N_5728[85]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [85])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1110.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1111 (.D(key_mem_0__127__N_5728[86]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [86])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1111.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1112 (.D(key_mem_0__127__N_5728[87]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [87])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1112.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1113 (.D(key_mem_0__127__N_5728[88]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [88])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1113.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1114 (.D(key_mem_0__127__N_5728[89]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [89])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1114.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1115 (.D(key_mem_0__127__N_5728[90]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [90])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1115.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1116 (.D(key_mem_0__127__N_5728[91]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [91])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1116.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1117 (.D(key_mem_0__127__N_5728[92]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [92])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1117.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1118 (.D(key_mem_0__127__N_5728[93]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [93])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1118.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1119 (.D(key_mem_0__127__N_5728[94]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [94])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1119.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1120 (.D(key_mem_0__127__N_5728[95]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [95])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1120.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1121 (.D(key_mem_0__127__N_5728[96]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [96])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1121.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1122 (.D(key_mem_0__127__N_5728[97]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [97])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1122.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1123 (.D(key_mem_0__127__N_5728[98]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [98])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1123.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1124 (.D(key_mem_0__127__N_5728[99]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [99])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1124.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1125 (.D(key_mem_0__127__N_5728[100]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [100])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1125.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1126 (.D(key_mem_0__127__N_5728[101]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [101])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1126.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1127 (.D(key_mem_0__127__N_5728[102]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [102])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1127.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1128 (.D(key_mem_0__127__N_5728[103]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [103])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1128.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1129 (.D(key_mem_0__127__N_5728[104]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [104])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1129.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1130 (.D(key_mem_0__127__N_5728[105]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [105])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1130.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1131 (.D(key_mem_0__127__N_5728[106]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [106])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1131.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1132 (.D(key_mem_0__127__N_5728[107]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [107])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1132.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1133 (.D(key_mem_0__127__N_5728[108]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [108])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1133.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1134 (.D(key_mem_0__127__N_5728[109]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [109])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1134.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1135 (.D(key_mem_0__127__N_5728[110]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [110])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1135.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1136 (.D(key_mem_0__127__N_5728[111]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [111])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1136.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1137 (.D(key_mem_0__127__N_5728[112]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [112])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1137.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1138 (.D(key_mem_0__127__N_5728[113]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [113])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1138.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1139 (.D(key_mem_0__127__N_5728[114]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [114])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1139.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1140 (.D(key_mem_0__127__N_5728[115]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [115])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1140.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1141 (.D(key_mem_0__127__N_5728[116]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [116])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1141.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1142 (.D(key_mem_0__127__N_5728[117]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [117])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1142.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1143 (.D(key_mem_0__127__N_5728[118]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [118])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1143.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1144 (.D(key_mem_0__127__N_5728[119]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [119])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1144.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1145 (.D(key_mem_0__127__N_5728[120]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [120])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1145.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1146 (.D(key_mem_0__127__N_5728[121]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [121])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1146.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1147 (.D(key_mem_0__127__N_5728[122]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [122])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1147.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1148 (.D(key_mem_0__127__N_5728[123]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [123])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1148.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1149 (.D(key_mem_0__127__N_5728[124]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [124])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1149.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1150 (.D(key_mem_0__127__N_5728[125]), .SP(clk_c_enable_1536), 
            .CK(clk_c), .Q(\key_mem[6] [125])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1150.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1151 (.D(key_mem_0__127__N_5728[126]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[6] [126])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1151.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1152 (.D(key_mem_0__127__N_5728[127]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[6] [127])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1152.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1153 (.D(key_mem_0__127__N_5600[0]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1153.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1154 (.D(key_mem_0__127__N_5600[1]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [1])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1154.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1155 (.D(key_mem_0__127__N_5600[2]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [2])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1155.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1156 (.D(key_mem_0__127__N_5600[3]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [3])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1156.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1157 (.D(key_mem_0__127__N_5600[4]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [4])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1157.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1158 (.D(key_mem_0__127__N_5600[5]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [5])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1158.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1159 (.D(key_mem_0__127__N_5600[6]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [6])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1159.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1160 (.D(key_mem_0__127__N_5600[7]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [7])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1160.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1161 (.D(key_mem_0__127__N_5600[8]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [8])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1161.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1162 (.D(key_mem_0__127__N_5600[9]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [9])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1162.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1163 (.D(key_mem_0__127__N_5600[10]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [10])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1163.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1164 (.D(key_mem_0__127__N_5600[11]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [11])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1164.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1165 (.D(key_mem_0__127__N_5600[12]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [12])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1165.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1166 (.D(key_mem_0__127__N_5600[13]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [13])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1166.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1167 (.D(key_mem_0__127__N_5600[14]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [14])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1167.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1168 (.D(key_mem_0__127__N_5600[15]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [15])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1168.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1169 (.D(key_mem_0__127__N_5600[16]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [16])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1169.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1170 (.D(key_mem_0__127__N_5600[17]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [17])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1170.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1171 (.D(key_mem_0__127__N_5600[18]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [18])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1171.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1172 (.D(key_mem_0__127__N_5600[19]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [19])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1172.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1173 (.D(key_mem_0__127__N_5600[20]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [20])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1173.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1174 (.D(key_mem_0__127__N_5600[21]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [21])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1174.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1175 (.D(key_mem_0__127__N_5600[22]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [22])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1175.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1176 (.D(key_mem_0__127__N_5600[23]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [23])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1176.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1177 (.D(key_mem_0__127__N_5600[24]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [24])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1177.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1178 (.D(key_mem_0__127__N_5600[25]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [25])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1178.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1179 (.D(key_mem_0__127__N_5600[26]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [26])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1179.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1180 (.D(key_mem_0__127__N_5600[27]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [27])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1180.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1181 (.D(key_mem_0__127__N_5600[28]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [28])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1181.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1182 (.D(key_mem_0__127__N_5600[29]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [29])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1182.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1183 (.D(key_mem_0__127__N_5600[30]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [30])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1183.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1184 (.D(key_mem_0__127__N_5600[31]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [31])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1184.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1185 (.D(key_mem_0__127__N_5600[32]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [32])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1185.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1186 (.D(key_mem_0__127__N_5600[33]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [33])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1186.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1187 (.D(key_mem_0__127__N_5600[34]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [34])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1187.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1188 (.D(key_mem_0__127__N_5600[35]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [35])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1188.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1189 (.D(key_mem_0__127__N_5600[36]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [36])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1189.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1190 (.D(key_mem_0__127__N_5600[37]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [37])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1190.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1191 (.D(key_mem_0__127__N_5600[38]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [38])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1191.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1192 (.D(key_mem_0__127__N_5600[39]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [39])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1192.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1193 (.D(key_mem_0__127__N_5600[40]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [40])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1193.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1194 (.D(key_mem_0__127__N_5600[41]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [41])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1194.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1195 (.D(key_mem_0__127__N_5600[42]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [42])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1195.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1196 (.D(key_mem_0__127__N_5600[43]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [43])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1196.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1197 (.D(key_mem_0__127__N_5600[44]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [44])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1197.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1198 (.D(key_mem_0__127__N_5600[45]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [45])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1198.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1199 (.D(key_mem_0__127__N_5600[46]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [46])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1199.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1200 (.D(key_mem_0__127__N_5600[47]), .SP(clk_c_enable_1586), 
            .CK(clk_c), .Q(\key_mem[5] [47])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1200.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1201 (.D(key_mem_0__127__N_5600[48]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [48])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1201.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1202 (.D(key_mem_0__127__N_5600[49]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [49])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1202.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1203 (.D(key_mem_0__127__N_5600[50]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [50])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1203.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1204 (.D(key_mem_0__127__N_5600[51]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [51])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1204.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1205 (.D(key_mem_0__127__N_5600[52]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [52])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1205.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1206 (.D(key_mem_0__127__N_5600[53]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [53])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1206.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1207 (.D(key_mem_0__127__N_5600[54]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [54])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1207.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1208 (.D(key_mem_0__127__N_5600[55]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [55])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1208.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1209 (.D(key_mem_0__127__N_5600[56]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [56])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1209.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1210 (.D(key_mem_0__127__N_5600[57]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [57])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1210.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1211 (.D(key_mem_0__127__N_5600[58]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [58])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1211.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1212 (.D(key_mem_0__127__N_5600[59]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [59])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1212.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1213 (.D(key_mem_0__127__N_5600[60]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [60])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1213.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1214 (.D(key_mem_0__127__N_5600[61]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [61])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1214.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1215 (.D(key_mem_0__127__N_5600[62]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [62])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1215.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1216 (.D(key_mem_0__127__N_5600[63]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [63])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1216.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1217 (.D(key_mem_0__127__N_5600[64]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [64])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1217.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1218 (.D(key_mem_0__127__N_5600[65]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [65])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1218.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1219 (.D(key_mem_0__127__N_5600[66]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [66])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1219.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1220 (.D(key_mem_0__127__N_5600[67]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [67])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1220.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1221 (.D(key_mem_0__127__N_5600[68]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [68])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1221.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1222 (.D(key_mem_0__127__N_5600[69]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [69])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1222.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1223 (.D(key_mem_0__127__N_5600[70]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [70])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1223.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1224 (.D(key_mem_0__127__N_5600[71]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [71])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1224.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1225 (.D(key_mem_0__127__N_5600[72]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [72])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1225.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1226 (.D(key_mem_0__127__N_5600[73]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [73])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1226.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1227 (.D(key_mem_0__127__N_5600[74]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [74])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1227.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1228 (.D(key_mem_0__127__N_5600[75]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [75])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1228.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1229 (.D(key_mem_0__127__N_5600[76]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [76])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1229.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1230 (.D(key_mem_0__127__N_5600[77]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [77])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1230.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1231 (.D(key_mem_0__127__N_5600[78]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [78])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1231.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1232 (.D(key_mem_0__127__N_5600[79]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [79])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1232.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1233 (.D(key_mem_0__127__N_5600[80]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [80])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1233.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1234 (.D(key_mem_0__127__N_5600[81]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [81])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1234.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1235 (.D(key_mem_0__127__N_5600[82]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [82])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1235.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1236 (.D(key_mem_0__127__N_5600[83]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [83])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1236.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1237 (.D(key_mem_0__127__N_5600[84]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [84])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1237.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1238 (.D(key_mem_0__127__N_5600[85]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [85])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1238.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1239 (.D(key_mem_0__127__N_5600[86]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [86])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1239.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1240 (.D(key_mem_0__127__N_5600[87]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [87])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1240.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1241 (.D(key_mem_0__127__N_5600[88]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [88])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1241.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1242 (.D(key_mem_0__127__N_5600[89]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [89])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1242.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1243 (.D(key_mem_0__127__N_5600[90]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [90])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1243.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1244 (.D(key_mem_0__127__N_5600[91]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [91])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1244.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1245 (.D(key_mem_0__127__N_5600[92]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [92])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1245.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1246 (.D(key_mem_0__127__N_5600[93]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [93])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1246.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1247 (.D(key_mem_0__127__N_5600[94]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [94])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1247.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1248 (.D(key_mem_0__127__N_5600[95]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [95])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1248.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1249 (.D(key_mem_0__127__N_5600[96]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [96])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1249.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1250 (.D(key_mem_0__127__N_5600[97]), .SP(clk_c_enable_1636), 
            .CK(clk_c), .Q(\key_mem[5] [97])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1250.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1251 (.D(key_mem_0__127__N_5600[98]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[5] [98])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1251.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1252 (.D(key_mem_0__127__N_5600[99]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[5] [99])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1252.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1253 (.D(key_mem_0__127__N_5600[100]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[5] [100])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1253.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1254 (.D(key_mem_0__127__N_5600[101]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[5] [101])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1254.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1255 (.D(key_mem_0__127__N_5600[102]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[5] [102])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1255.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1256 (.D(key_mem_0__127__N_5600[103]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[5] [103])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1256.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1257 (.D(key_mem_0__127__N_5600[104]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[5] [104])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1257.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1258 (.D(key_mem_0__127__N_5600[105]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[5] [105])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1258.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1259 (.D(key_mem_0__127__N_5600[106]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[5] [106])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1259.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1260 (.D(key_mem_0__127__N_5600[107]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[5] [107])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1260.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1261 (.D(key_mem_0__127__N_5600[108]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[5] [108])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1261.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1262 (.D(key_mem_0__127__N_5600[109]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[5] [109])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1262.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1263 (.D(key_mem_0__127__N_5600[110]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[5] [110])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1263.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1264 (.D(key_mem_0__127__N_5600[111]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[5] [111])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1264.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1265 (.D(key_mem_0__127__N_5600[112]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[5] [112])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1265.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1266 (.D(key_mem_0__127__N_5600[113]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[5] [113])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1266.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1267 (.D(key_mem_0__127__N_5600[114]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[5] [114])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1267.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1268 (.D(key_mem_0__127__N_5600[115]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[5] [115])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1268.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1269 (.D(key_mem_0__127__N_5600[116]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[5] [116])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1269.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1270 (.D(key_mem_0__127__N_5600[117]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[5] [117])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1270.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1271 (.D(key_mem_0__127__N_5600[118]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[5] [118])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1271.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1272 (.D(key_mem_0__127__N_5600[119]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[5] [119])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1272.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1273 (.D(key_mem_0__127__N_5600[120]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[5] [120])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1273.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1274 (.D(key_mem_0__127__N_5600[121]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[5] [121])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1274.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1275 (.D(key_mem_0__127__N_5600[122]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[5] [122])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1275.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1276 (.D(key_mem_0__127__N_5600[123]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[5] [123])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1276.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1277 (.D(key_mem_0__127__N_5600[124]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[5] [124])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1277.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1278 (.D(key_mem_0__127__N_5600[125]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[5] [125])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1278.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1279 (.D(key_mem_0__127__N_5600[126]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[5] [126])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1279.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1280 (.D(key_mem_0__127__N_5600[127]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[5] [127])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1280.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1281 (.D(key_mem_0__127__N_5472[0]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[4] [0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1281.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1282 (.D(key_mem_0__127__N_5472[1]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[4] [1])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1282.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1283 (.D(key_mem_0__127__N_5472[2]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[4] [2])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1283.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1284 (.D(key_mem_0__127__N_5472[3]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[4] [3])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1284.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1285 (.D(key_mem_0__127__N_5472[4]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[4] [4])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1285.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1286 (.D(key_mem_0__127__N_5472[5]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[4] [5])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1286.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1287 (.D(key_mem_0__127__N_5472[6]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[4] [6])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1287.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1288 (.D(key_mem_0__127__N_5472[7]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[4] [7])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1288.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1289 (.D(key_mem_0__127__N_5472[8]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[4] [8])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1289.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1290 (.D(key_mem_0__127__N_5472[9]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[4] [9])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1290.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1291 (.D(key_mem_0__127__N_5472[10]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[4] [10])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1291.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1292 (.D(key_mem_0__127__N_5472[11]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[4] [11])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1292.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1293 (.D(key_mem_0__127__N_5472[12]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[4] [12])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1293.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1294 (.D(key_mem_0__127__N_5472[13]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[4] [13])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1294.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1295 (.D(key_mem_0__127__N_5472[14]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[4] [14])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1295.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1296 (.D(key_mem_0__127__N_5472[15]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[4] [15])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1296.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1297 (.D(key_mem_0__127__N_5472[16]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[4] [16])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1297.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1298 (.D(key_mem_0__127__N_5472[17]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[4] [17])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1298.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1299 (.D(key_mem_0__127__N_5472[18]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[4] [18])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1299.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1300 (.D(key_mem_0__127__N_5472[19]), .SP(clk_c_enable_1686), 
            .CK(clk_c), .Q(\key_mem[4] [19])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1300.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1301 (.D(key_mem_0__127__N_5472[20]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [20])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1301.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1302 (.D(key_mem_0__127__N_5472[21]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [21])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1302.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1303 (.D(key_mem_0__127__N_5472[22]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [22])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1303.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1304 (.D(key_mem_0__127__N_5472[23]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [23])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1304.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1305 (.D(key_mem_0__127__N_5472[24]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [24])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1305.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1306 (.D(key_mem_0__127__N_5472[25]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [25])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1306.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1307 (.D(key_mem_0__127__N_5472[26]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [26])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1307.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1308 (.D(key_mem_0__127__N_5472[27]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [27])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1308.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1309 (.D(key_mem_0__127__N_5472[28]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [28])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1309.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1310 (.D(key_mem_0__127__N_5472[29]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [29])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1310.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1311 (.D(key_mem_0__127__N_5472[30]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [30])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1311.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1312 (.D(key_mem_0__127__N_5472[31]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [31])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1312.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1313 (.D(key_mem_0__127__N_5472[32]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [32])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1313.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1314 (.D(key_mem_0__127__N_5472[33]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [33])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1314.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1315 (.D(key_mem_0__127__N_5472[34]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [34])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1315.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1316 (.D(key_mem_0__127__N_5472[35]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [35])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1316.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1317 (.D(key_mem_0__127__N_5472[36]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [36])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1317.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1318 (.D(key_mem_0__127__N_5472[37]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [37])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1318.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1319 (.D(key_mem_0__127__N_5472[38]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [38])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1319.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1320 (.D(key_mem_0__127__N_5472[39]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [39])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1320.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1321 (.D(key_mem_0__127__N_5472[40]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [40])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1321.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1322 (.D(key_mem_0__127__N_5472[41]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [41])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1322.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1323 (.D(key_mem_0__127__N_5472[42]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [42])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1323.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1324 (.D(key_mem_0__127__N_5472[43]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [43])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1324.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1325 (.D(key_mem_0__127__N_5472[44]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [44])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1325.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1326 (.D(key_mem_0__127__N_5472[45]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [45])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1326.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1327 (.D(key_mem_0__127__N_5472[46]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [46])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1327.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1328 (.D(key_mem_0__127__N_5472[47]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [47])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1328.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1329 (.D(key_mem_0__127__N_5472[48]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [48])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1329.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1330 (.D(key_mem_0__127__N_5472[49]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [49])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1330.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1331 (.D(key_mem_0__127__N_5472[50]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [50])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1331.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1332 (.D(key_mem_0__127__N_5472[51]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [51])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1332.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1333 (.D(key_mem_0__127__N_5472[52]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [52])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1333.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1334 (.D(key_mem_0__127__N_5472[53]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [53])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1334.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1335 (.D(key_mem_0__127__N_5472[54]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [54])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1335.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1336 (.D(key_mem_0__127__N_5472[55]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [55])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1336.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1337 (.D(key_mem_0__127__N_5472[56]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [56])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1337.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1338 (.D(key_mem_0__127__N_5472[57]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [57])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1338.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1339 (.D(key_mem_0__127__N_5472[58]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [58])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1339.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1340 (.D(key_mem_0__127__N_5472[59]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [59])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1340.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1341 (.D(key_mem_0__127__N_5472[60]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [60])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1341.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1342 (.D(key_mem_0__127__N_5472[61]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [61])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1342.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1343 (.D(key_mem_0__127__N_5472[62]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [62])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1343.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1344 (.D(key_mem_0__127__N_5472[63]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [63])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1344.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1345 (.D(key_mem_0__127__N_5472[64]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [64])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1345.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1346 (.D(key_mem_0__127__N_5472[65]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [65])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1346.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1347 (.D(key_mem_0__127__N_5472[66]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [66])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1347.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1348 (.D(key_mem_0__127__N_5472[67]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [67])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1348.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1349 (.D(key_mem_0__127__N_5472[68]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [68])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1349.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1350 (.D(key_mem_0__127__N_5472[69]), .SP(clk_c_enable_1736), 
            .CK(clk_c), .Q(\key_mem[4] [69])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1350.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1351 (.D(key_mem_0__127__N_5472[70]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [70])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1351.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1352 (.D(key_mem_0__127__N_5472[71]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [71])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1352.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1353 (.D(key_mem_0__127__N_5472[72]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [72])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1353.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1354 (.D(key_mem_0__127__N_5472[73]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [73])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1354.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1355 (.D(key_mem_0__127__N_5472[74]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [74])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1355.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1356 (.D(key_mem_0__127__N_5472[75]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [75])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1356.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1357 (.D(key_mem_0__127__N_5472[76]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [76])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1357.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1358 (.D(key_mem_0__127__N_5472[77]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [77])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1358.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1359 (.D(key_mem_0__127__N_5472[78]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [78])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1359.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1360 (.D(key_mem_0__127__N_5472[79]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [79])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1360.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1361 (.D(key_mem_0__127__N_5472[80]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [80])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1361.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1362 (.D(key_mem_0__127__N_5472[81]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [81])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1362.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1363 (.D(key_mem_0__127__N_5472[82]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [82])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1363.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1364 (.D(key_mem_0__127__N_5472[83]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [83])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1364.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1365 (.D(key_mem_0__127__N_5472[84]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [84])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1365.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1366 (.D(key_mem_0__127__N_5472[85]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [85])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1366.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1367 (.D(key_mem_0__127__N_5472[86]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [86])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1367.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1368 (.D(key_mem_0__127__N_5472[87]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [87])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1368.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1369 (.D(key_mem_0__127__N_5472[88]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [88])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1369.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1370 (.D(key_mem_0__127__N_5472[89]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [89])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1370.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1371 (.D(key_mem_0__127__N_5472[90]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [90])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1371.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1372 (.D(key_mem_0__127__N_5472[91]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [91])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1372.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1373 (.D(key_mem_0__127__N_5472[92]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [92])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1373.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1374 (.D(key_mem_0__127__N_5472[93]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [93])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1374.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1375 (.D(key_mem_0__127__N_5472[94]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [94])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1375.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1376 (.D(key_mem_0__127__N_5472[95]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [95])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1376.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1377 (.D(key_mem_0__127__N_5472[96]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [96])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1377.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1378 (.D(key_mem_0__127__N_5472[97]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [97])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1378.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1379 (.D(key_mem_0__127__N_5472[98]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [98])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1379.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1380 (.D(key_mem_0__127__N_5472[99]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [99])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1380.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1381 (.D(key_mem_0__127__N_5472[100]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [100])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1381.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1382 (.D(key_mem_0__127__N_5472[101]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [101])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1382.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1383 (.D(key_mem_0__127__N_5472[102]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [102])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1383.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1384 (.D(key_mem_0__127__N_5472[103]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [103])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1384.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1385 (.D(key_mem_0__127__N_5472[104]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [104])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1385.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1386 (.D(key_mem_0__127__N_5472[105]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [105])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1386.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1387 (.D(key_mem_0__127__N_5472[106]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [106])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1387.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1388 (.D(key_mem_0__127__N_5472[107]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [107])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1388.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1389 (.D(key_mem_0__127__N_5472[108]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [108])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1389.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1390 (.D(key_mem_0__127__N_5472[109]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [109])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1390.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1391 (.D(key_mem_0__127__N_5472[110]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [110])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1391.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1392 (.D(key_mem_0__127__N_5472[111]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [111])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1392.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1393 (.D(key_mem_0__127__N_5472[112]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [112])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1393.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1394 (.D(key_mem_0__127__N_5472[113]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [113])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1394.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1395 (.D(key_mem_0__127__N_5472[114]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [114])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1395.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1396 (.D(key_mem_0__127__N_5472[115]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [115])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1396.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1397 (.D(key_mem_0__127__N_5472[116]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [116])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1397.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1398 (.D(key_mem_0__127__N_5472[117]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [117])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1398.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1399 (.D(key_mem_0__127__N_5472[118]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [118])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1399.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1400 (.D(key_mem_0__127__N_5472[119]), .SP(clk_c_enable_1786), 
            .CK(clk_c), .Q(\key_mem[4] [119])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1400.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1401 (.D(key_mem_0__127__N_5472[120]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[4] [120])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1401.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1402 (.D(key_mem_0__127__N_5472[121]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[4] [121])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1402.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1403 (.D(key_mem_0__127__N_5472[122]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[4] [122])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1403.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1404 (.D(key_mem_0__127__N_5472[123]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[4] [123])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1404.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1405 (.D(key_mem_0__127__N_5472[124]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[4] [124])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1405.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1406 (.D(key_mem_0__127__N_5472[125]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[4] [125])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1406.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1407 (.D(key_mem_0__127__N_5472[126]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[4] [126])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1407.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1408 (.D(key_mem_0__127__N_5472[127]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[4] [127])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1408.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1409 (.D(key_mem_0__127__N_5344[0]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[3] [0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1409.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1410 (.D(key_mem_0__127__N_5344[1]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[3] [1])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1410.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1411 (.D(key_mem_0__127__N_5344[2]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[3] [2])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1411.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1412 (.D(key_mem_0__127__N_5344[3]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[3] [3])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1412.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1413 (.D(key_mem_0__127__N_5344[4]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[3] [4])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1413.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1414 (.D(key_mem_0__127__N_5344[5]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[3] [5])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1414.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1415 (.D(key_mem_0__127__N_5344[6]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[3] [6])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1415.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1416 (.D(key_mem_0__127__N_5344[7]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[3] [7])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1416.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1417 (.D(key_mem_0__127__N_5344[8]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[3] [8])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1417.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1418 (.D(key_mem_0__127__N_5344[9]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[3] [9])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1418.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1419 (.D(key_mem_0__127__N_5344[10]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[3] [10])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1419.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1420 (.D(key_mem_0__127__N_5344[11]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[3] [11])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1420.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1421 (.D(key_mem_0__127__N_5344[12]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[3] [12])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1421.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1422 (.D(key_mem_0__127__N_5344[13]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[3] [13])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1422.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1423 (.D(key_mem_0__127__N_5344[14]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[3] [14])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1423.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1424 (.D(key_mem_0__127__N_5344[15]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[3] [15])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1424.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1425 (.D(key_mem_0__127__N_5344[16]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[3] [16])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1425.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1426 (.D(key_mem_0__127__N_5344[17]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[3] [17])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1426.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1427 (.D(key_mem_0__127__N_5344[18]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[3] [18])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1427.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1428 (.D(key_mem_0__127__N_5344[19]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[3] [19])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1428.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1429 (.D(key_mem_0__127__N_5344[20]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[3] [20])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1429.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1430 (.D(key_mem_0__127__N_5344[21]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[3] [21])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1430.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1431 (.D(key_mem_0__127__N_5344[22]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[3] [22])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1431.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1432 (.D(key_mem_0__127__N_5344[23]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[3] [23])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1432.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1433 (.D(key_mem_0__127__N_5344[24]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[3] [24])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1433.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1434 (.D(key_mem_0__127__N_5344[25]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[3] [25])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1434.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1435 (.D(key_mem_0__127__N_5344[26]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[3] [26])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1435.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1436 (.D(key_mem_0__127__N_5344[27]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[3] [27])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1436.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1437 (.D(key_mem_0__127__N_5344[28]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[3] [28])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1437.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1438 (.D(key_mem_0__127__N_5344[29]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[3] [29])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1438.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1439 (.D(key_mem_0__127__N_5344[30]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[3] [30])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1439.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1440 (.D(key_mem_0__127__N_5344[31]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[3] [31])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1440.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1441 (.D(key_mem_0__127__N_5344[32]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[3] [32])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1441.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1442 (.D(key_mem_0__127__N_5344[33]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[3] [33])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1442.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1443 (.D(key_mem_0__127__N_5344[34]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[3] [34])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1443.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1444 (.D(key_mem_0__127__N_5344[35]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[3] [35])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1444.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1445 (.D(key_mem_0__127__N_5344[36]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[3] [36])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1445.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1446 (.D(key_mem_0__127__N_5344[37]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[3] [37])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1446.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1447 (.D(key_mem_0__127__N_5344[38]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[3] [38])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1447.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1448 (.D(key_mem_0__127__N_5344[39]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[3] [39])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1448.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1449 (.D(key_mem_0__127__N_5344[40]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[3] [40])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1449.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1450 (.D(key_mem_0__127__N_5344[41]), .SP(clk_c_enable_1836), 
            .CK(clk_c), .Q(\key_mem[3] [41])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1450.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1451 (.D(key_mem_0__127__N_5344[42]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [42])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1451.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1452 (.D(key_mem_0__127__N_5344[43]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [43])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1452.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1453 (.D(key_mem_0__127__N_5344[44]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [44])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1453.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1454 (.D(key_mem_0__127__N_5344[45]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [45])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1454.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1455 (.D(key_mem_0__127__N_5344[46]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [46])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1455.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1456 (.D(key_mem_0__127__N_5344[47]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [47])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1456.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1457 (.D(key_mem_0__127__N_5344[48]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [48])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1457.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1458 (.D(key_mem_0__127__N_5344[49]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [49])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1458.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1459 (.D(key_mem_0__127__N_5344[50]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [50])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1459.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1460 (.D(key_mem_0__127__N_5344[51]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [51])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1460.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1461 (.D(key_mem_0__127__N_5344[52]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [52])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1461.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1462 (.D(key_mem_0__127__N_5344[53]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [53])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1462.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1463 (.D(key_mem_0__127__N_5344[54]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [54])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1463.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1464 (.D(key_mem_0__127__N_5344[55]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [55])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1464.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1465 (.D(key_mem_0__127__N_5344[56]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [56])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1465.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1466 (.D(key_mem_0__127__N_5344[57]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [57])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1466.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1467 (.D(key_mem_0__127__N_5344[58]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [58])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1467.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1468 (.D(key_mem_0__127__N_5344[59]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [59])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1468.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1469 (.D(key_mem_0__127__N_5344[60]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [60])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1469.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1470 (.D(key_mem_0__127__N_5344[61]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [61])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1470.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1471 (.D(key_mem_0__127__N_5344[62]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [62])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1471.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1472 (.D(key_mem_0__127__N_5344[63]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [63])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1472.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1473 (.D(key_mem_0__127__N_5344[64]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [64])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1473.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1474 (.D(key_mem_0__127__N_5344[65]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [65])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1474.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1475 (.D(key_mem_0__127__N_5344[66]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [66])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1475.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1476 (.D(key_mem_0__127__N_5344[67]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [67])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1476.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1477 (.D(key_mem_0__127__N_5344[68]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [68])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1477.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1478 (.D(key_mem_0__127__N_5344[69]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [69])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1478.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1479 (.D(key_mem_0__127__N_5344[70]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [70])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1479.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1480 (.D(key_mem_0__127__N_5344[71]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [71])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1480.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1481 (.D(key_mem_0__127__N_5344[72]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [72])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1481.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1482 (.D(key_mem_0__127__N_5344[73]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [73])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1482.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1483 (.D(key_mem_0__127__N_5344[74]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [74])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1483.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1484 (.D(key_mem_0__127__N_5344[75]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [75])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1484.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1485 (.D(key_mem_0__127__N_5344[76]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [76])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1485.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1486 (.D(key_mem_0__127__N_5344[77]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [77])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1486.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1487 (.D(key_mem_0__127__N_5344[78]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [78])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1487.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1488 (.D(key_mem_0__127__N_5344[79]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [79])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1488.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1489 (.D(key_mem_0__127__N_5344[80]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [80])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1489.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1490 (.D(key_mem_0__127__N_5344[81]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [81])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1490.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1491 (.D(key_mem_0__127__N_5344[82]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [82])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1491.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1492 (.D(key_mem_0__127__N_5344[83]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [83])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1492.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1493 (.D(key_mem_0__127__N_5344[84]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [84])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1493.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1494 (.D(key_mem_0__127__N_5344[85]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [85])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1494.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1495 (.D(key_mem_0__127__N_5344[86]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [86])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1495.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1496 (.D(key_mem_0__127__N_5344[87]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [87])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1496.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1497 (.D(key_mem_0__127__N_5344[88]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [88])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1497.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1498 (.D(key_mem_0__127__N_5344[89]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [89])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1498.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1499 (.D(key_mem_0__127__N_5344[90]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [90])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1499.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1500 (.D(key_mem_0__127__N_5344[91]), .SP(clk_c_enable_1886), 
            .CK(clk_c), .Q(\key_mem[3] [91])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1500.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1501 (.D(key_mem_0__127__N_5344[92]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[3] [92])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1501.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1502 (.D(key_mem_0__127__N_5344[93]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[3] [93])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1502.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1503 (.D(key_mem_0__127__N_5344[94]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[3] [94])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1503.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1504 (.D(key_mem_0__127__N_5344[95]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[3] [95])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1504.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1505 (.D(key_mem_0__127__N_5344[96]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[3] [96])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1505.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1506 (.D(key_mem_0__127__N_5344[97]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[3] [97])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1506.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1507 (.D(key_mem_0__127__N_5344[98]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[3] [98])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1507.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1508 (.D(key_mem_0__127__N_5344[99]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[3] [99])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1508.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1509 (.D(key_mem_0__127__N_5344[100]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[3] [100])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1509.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1510 (.D(key_mem_0__127__N_5344[101]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[3] [101])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1510.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1511 (.D(key_mem_0__127__N_5344[102]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[3] [102])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1511.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1512 (.D(key_mem_0__127__N_5344[103]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[3] [103])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1512.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1513 (.D(key_mem_0__127__N_5344[104]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[3] [104])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1513.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1514 (.D(key_mem_0__127__N_5344[105]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[3] [105])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1514.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1515 (.D(key_mem_0__127__N_5344[106]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[3] [106])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1515.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1516 (.D(key_mem_0__127__N_5344[107]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[3] [107])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1516.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1517 (.D(key_mem_0__127__N_5344[108]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[3] [108])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1517.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1518 (.D(key_mem_0__127__N_5344[109]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[3] [109])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1518.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1519 (.D(key_mem_0__127__N_5344[110]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[3] [110])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1519.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1520 (.D(key_mem_0__127__N_5344[111]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[3] [111])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1520.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1521 (.D(key_mem_0__127__N_5344[112]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[3] [112])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1521.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1522 (.D(key_mem_0__127__N_5344[113]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[3] [113])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1522.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1523 (.D(key_mem_0__127__N_5344[114]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[3] [114])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1523.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1524 (.D(key_mem_0__127__N_5344[115]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[3] [115])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1524.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1525 (.D(key_mem_0__127__N_5344[116]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[3] [116])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1525.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1526 (.D(key_mem_0__127__N_5344[117]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[3] [117])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1526.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1527 (.D(key_mem_0__127__N_5344[118]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[3] [118])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1527.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1528 (.D(key_mem_0__127__N_5344[119]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[3] [119])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1528.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1529 (.D(key_mem_0__127__N_5344[120]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[3] [120])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1529.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1530 (.D(key_mem_0__127__N_5344[121]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[3] [121])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1530.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1531 (.D(key_mem_0__127__N_5344[122]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[3] [122])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1531.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1532 (.D(key_mem_0__127__N_5344[123]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[3] [123])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1532.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1533 (.D(key_mem_0__127__N_5344[124]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[3] [124])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1533.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1534 (.D(key_mem_0__127__N_5344[125]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[3] [125])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1534.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1535 (.D(key_mem_0__127__N_5344[126]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[3] [126])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1535.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1536 (.D(key_mem_0__127__N_5344[127]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[3] [127])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1536.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1537 (.D(key_mem_0__127__N_5216[0]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[2] [0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1537.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1538 (.D(key_mem_0__127__N_5216[1]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[2] [1])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1538.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1539 (.D(key_mem_0__127__N_5216[2]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[2] [2])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1539.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1540 (.D(key_mem_0__127__N_5216[3]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[2] [3])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1540.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1541 (.D(key_mem_0__127__N_5216[4]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[2] [4])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1541.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1542 (.D(key_mem_0__127__N_5216[5]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[2] [5])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1542.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1543 (.D(key_mem_0__127__N_5216[6]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[2] [6])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1543.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1544 (.D(key_mem_0__127__N_5216[7]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[2] [7])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1544.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1545 (.D(key_mem_0__127__N_5216[8]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[2] [8])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1545.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1546 (.D(key_mem_0__127__N_5216[9]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[2] [9])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1546.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1547 (.D(key_mem_0__127__N_5216[10]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[2] [10])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1547.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1548 (.D(key_mem_0__127__N_5216[11]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[2] [11])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1548.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1549 (.D(key_mem_0__127__N_5216[12]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[2] [12])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1549.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1550 (.D(key_mem_0__127__N_5216[13]), .SP(clk_c_enable_1936), 
            .CK(clk_c), .Q(\key_mem[2] [13])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1550.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1551 (.D(key_mem_0__127__N_5216[14]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [14])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1551.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1552 (.D(key_mem_0__127__N_5216[15]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [15])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1552.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1553 (.D(key_mem_0__127__N_5216[16]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [16])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1553.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1554 (.D(key_mem_0__127__N_5216[17]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [17])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1554.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1555 (.D(key_mem_0__127__N_5216[18]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [18])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1555.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1556 (.D(key_mem_0__127__N_5216[19]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [19])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1556.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1557 (.D(key_mem_0__127__N_5216[20]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [20])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1557.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1558 (.D(key_mem_0__127__N_5216[21]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [21])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1558.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1559 (.D(key_mem_0__127__N_5216[22]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [22])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1559.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1560 (.D(key_mem_0__127__N_5216[23]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [23])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1560.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1561 (.D(key_mem_0__127__N_5216[24]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [24])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1561.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1562 (.D(key_mem_0__127__N_5216[25]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [25])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1562.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1563 (.D(key_mem_0__127__N_5216[26]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [26])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1563.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1564 (.D(key_mem_0__127__N_5216[27]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [27])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1564.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1565 (.D(key_mem_0__127__N_5216[28]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [28])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1565.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1566 (.D(key_mem_0__127__N_5216[29]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [29])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1566.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1567 (.D(key_mem_0__127__N_5216[30]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [30])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1567.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1568 (.D(key_mem_0__127__N_5216[31]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [31])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1568.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1569 (.D(key_mem_0__127__N_5216[32]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [32])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1569.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1570 (.D(key_mem_0__127__N_5216[33]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [33])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1570.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1571 (.D(key_mem_0__127__N_5216[34]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [34])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1571.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1572 (.D(key_mem_0__127__N_5216[35]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [35])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1572.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1573 (.D(key_mem_0__127__N_5216[36]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [36])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1573.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1574 (.D(key_mem_0__127__N_5216[37]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [37])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1574.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1575 (.D(key_mem_0__127__N_5216[38]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [38])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1575.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1576 (.D(key_mem_0__127__N_5216[39]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [39])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1576.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1577 (.D(key_mem_0__127__N_5216[40]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [40])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1577.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1578 (.D(key_mem_0__127__N_5216[41]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [41])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1578.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1579 (.D(key_mem_0__127__N_5216[42]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [42])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1579.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1580 (.D(key_mem_0__127__N_5216[43]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [43])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1580.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1581 (.D(key_mem_0__127__N_5216[44]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [44])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1581.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1582 (.D(key_mem_0__127__N_5216[45]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [45])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1582.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1583 (.D(key_mem_0__127__N_5216[46]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [46])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1583.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1584 (.D(key_mem_0__127__N_5216[47]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [47])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1584.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1585 (.D(key_mem_0__127__N_5216[48]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [48])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1585.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1586 (.D(key_mem_0__127__N_5216[49]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [49])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1586.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1587 (.D(key_mem_0__127__N_5216[50]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [50])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1587.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1588 (.D(key_mem_0__127__N_5216[51]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [51])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1588.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1589 (.D(key_mem_0__127__N_5216[52]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [52])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1589.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1590 (.D(key_mem_0__127__N_5216[53]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [53])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1590.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1591 (.D(key_mem_0__127__N_5216[54]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [54])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1591.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1592 (.D(key_mem_0__127__N_5216[55]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [55])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1592.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1593 (.D(key_mem_0__127__N_5216[56]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [56])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1593.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1594 (.D(key_mem_0__127__N_5216[57]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [57])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1594.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1595 (.D(key_mem_0__127__N_5216[58]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [58])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1595.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1596 (.D(key_mem_0__127__N_5216[59]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [59])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1596.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1597 (.D(key_mem_0__127__N_5216[60]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [60])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1597.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1598 (.D(key_mem_0__127__N_5216[61]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [61])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1598.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1599 (.D(key_mem_0__127__N_5216[62]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [62])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1599.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1600 (.D(key_mem_0__127__N_5216[63]), .SP(clk_c_enable_1986), 
            .CK(clk_c), .Q(\key_mem[2] [63])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1600.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1601 (.D(key_mem_0__127__N_5216[64]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [64])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1601.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1602 (.D(key_mem_0__127__N_5216[65]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [65])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1602.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1603 (.D(key_mem_0__127__N_5216[66]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [66])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1603.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1604 (.D(key_mem_0__127__N_5216[67]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [67])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1604.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1605 (.D(key_mem_0__127__N_5216[68]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [68])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1605.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1606 (.D(key_mem_0__127__N_5216[69]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [69])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1606.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1607 (.D(key_mem_0__127__N_5216[70]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [70])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1607.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1608 (.D(key_mem_0__127__N_5216[71]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [71])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1608.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1609 (.D(key_mem_0__127__N_5216[72]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [72])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1609.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1610 (.D(key_mem_0__127__N_5216[73]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [73])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1610.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1611 (.D(key_mem_0__127__N_5216[74]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [74])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1611.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1612 (.D(key_mem_0__127__N_5216[75]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [75])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1612.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1613 (.D(key_mem_0__127__N_5216[76]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [76])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1613.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1614 (.D(key_mem_0__127__N_5216[77]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [77])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1614.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1615 (.D(key_mem_0__127__N_5216[78]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [78])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1615.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1616 (.D(key_mem_0__127__N_5216[79]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [79])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1616.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1617 (.D(key_mem_0__127__N_5216[80]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [80])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1617.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1618 (.D(key_mem_0__127__N_5216[81]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [81])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1618.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1619 (.D(key_mem_0__127__N_5216[82]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [82])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1619.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1620 (.D(key_mem_0__127__N_5216[83]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [83])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1620.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1621 (.D(key_mem_0__127__N_5216[84]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [84])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1621.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1622 (.D(key_mem_0__127__N_5216[85]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [85])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1622.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1623 (.D(key_mem_0__127__N_5216[86]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [86])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1623.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1624 (.D(key_mem_0__127__N_5216[87]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [87])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1624.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1625 (.D(key_mem_0__127__N_5216[88]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [88])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1625.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1626 (.D(key_mem_0__127__N_5216[89]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [89])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1626.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1627 (.D(key_mem_0__127__N_5216[90]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [90])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1627.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1628 (.D(key_mem_0__127__N_5216[91]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [91])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1628.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1629 (.D(key_mem_0__127__N_5216[92]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [92])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1629.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1630 (.D(key_mem_0__127__N_5216[93]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [93])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1630.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1631 (.D(key_mem_0__127__N_5216[94]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [94])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1631.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1632 (.D(key_mem_0__127__N_5216[95]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [95])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1632.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1633 (.D(key_mem_0__127__N_5216[96]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [96])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1633.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1634 (.D(key_mem_0__127__N_5216[97]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [97])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1634.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1635 (.D(key_mem_0__127__N_5216[98]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [98])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1635.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1636 (.D(key_mem_0__127__N_5216[99]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [99])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1636.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1637 (.D(key_mem_0__127__N_5216[100]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [100])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1637.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1638 (.D(key_mem_0__127__N_5216[101]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [101])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1638.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1639 (.D(key_mem_0__127__N_5216[102]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [102])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1639.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1640 (.D(key_mem_0__127__N_5216[103]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [103])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1640.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1641 (.D(key_mem_0__127__N_5216[104]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [104])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1641.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1642 (.D(key_mem_0__127__N_5216[105]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [105])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1642.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1643 (.D(key_mem_0__127__N_5216[106]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [106])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1643.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1644 (.D(key_mem_0__127__N_5216[107]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [107])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1644.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1645 (.D(key_mem_0__127__N_5216[108]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [108])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1645.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1646 (.D(key_mem_0__127__N_5216[109]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [109])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1646.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1647 (.D(key_mem_0__127__N_5216[110]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [110])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1647.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1648 (.D(key_mem_0__127__N_5216[111]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [111])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1648.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1649 (.D(key_mem_0__127__N_5216[112]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [112])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1649.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1650 (.D(key_mem_0__127__N_5216[113]), .SP(clk_c_enable_2036), 
            .CK(clk_c), .Q(\key_mem[2] [113])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1650.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1651 (.D(key_mem_0__127__N_5216[114]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[2] [114])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1651.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1652 (.D(key_mem_0__127__N_5216[115]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[2] [115])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1652.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1653 (.D(key_mem_0__127__N_5216[116]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[2] [116])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1653.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1654 (.D(key_mem_0__127__N_5216[117]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[2] [117])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1654.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1655 (.D(key_mem_0__127__N_5216[118]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[2] [118])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1655.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1656 (.D(key_mem_0__127__N_5216[119]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[2] [119])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1656.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1657 (.D(key_mem_0__127__N_5216[120]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[2] [120])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1657.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1658 (.D(key_mem_0__127__N_5216[121]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[2] [121])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1658.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1659 (.D(key_mem_0__127__N_5216[122]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[2] [122])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1659.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1660 (.D(key_mem_0__127__N_5216[123]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[2] [123])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1660.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1661 (.D(key_mem_0__127__N_5216[124]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[2] [124])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1661.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1662 (.D(key_mem_0__127__N_5216[125]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[2] [125])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1662.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1663 (.D(key_mem_0__127__N_5216[126]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[2] [126])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1663.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1664 (.D(key_mem_0__127__N_5216[127]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[2] [127])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1664.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1665 (.D(key_mem_0__127__N_5088[0]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[1] [0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1665.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1666 (.D(key_mem_0__127__N_5088[1]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[1] [1])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1666.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1667 (.D(key_mem_0__127__N_5088[2]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[1] [2])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1667.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1668 (.D(key_mem_0__127__N_5088[3]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[1] [3])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1668.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1669 (.D(key_mem_0__127__N_5088[4]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[1] [4])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1669.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1670 (.D(key_mem_0__127__N_5088[5]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[1] [5])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1670.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1671 (.D(key_mem_0__127__N_5088[6]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[1] [6])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1671.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1672 (.D(key_mem_0__127__N_5088[7]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[1] [7])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1672.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1673 (.D(key_mem_0__127__N_5088[8]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[1] [8])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1673.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1674 (.D(key_mem_0__127__N_5088[9]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[1] [9])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1674.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1675 (.D(key_mem_0__127__N_5088[10]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[1] [10])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1675.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1676 (.D(key_mem_0__127__N_5088[11]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[1] [11])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1676.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1677 (.D(key_mem_0__127__N_5088[12]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[1] [12])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1677.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1678 (.D(key_mem_0__127__N_5088[13]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[1] [13])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1678.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1679 (.D(key_mem_0__127__N_5088[14]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[1] [14])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1679.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1680 (.D(key_mem_0__127__N_5088[15]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[1] [15])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1680.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1681 (.D(key_mem_0__127__N_5088[16]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[1] [16])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1681.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1682 (.D(key_mem_0__127__N_5088[17]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[1] [17])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1682.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1683 (.D(key_mem_0__127__N_5088[18]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[1] [18])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1683.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1684 (.D(key_mem_0__127__N_5088[19]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[1] [19])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1684.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1685 (.D(key_mem_0__127__N_5088[20]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[1] [20])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1685.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1686 (.D(key_mem_0__127__N_5088[21]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[1] [21])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1686.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1687 (.D(key_mem_0__127__N_5088[22]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[1] [22])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1687.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1688 (.D(key_mem_0__127__N_5088[23]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[1] [23])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1688.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1689 (.D(key_mem_0__127__N_5088[24]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[1] [24])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1689.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1690 (.D(key_mem_0__127__N_5088[25]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[1] [25])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1690.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1691 (.D(key_mem_0__127__N_5088[26]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[1] [26])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1691.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1692 (.D(key_mem_0__127__N_5088[27]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[1] [27])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1692.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1693 (.D(key_mem_0__127__N_5088[28]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[1] [28])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1693.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1694 (.D(key_mem_0__127__N_5088[29]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[1] [29])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1694.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1695 (.D(key_mem_0__127__N_5088[30]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[1] [30])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1695.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1696 (.D(key_mem_0__127__N_5088[31]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[1] [31])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1696.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1697 (.D(key_mem_0__127__N_5088[32]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[1] [32])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1697.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1698 (.D(key_mem_0__127__N_5088[33]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[1] [33])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1698.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1699 (.D(key_mem_0__127__N_5088[34]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[1] [34])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1699.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1700 (.D(key_mem_0__127__N_5088[35]), .SP(clk_c_enable_2086), 
            .CK(clk_c), .Q(\key_mem[1] [35])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1700.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1701 (.D(key_mem_0__127__N_5088[36]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [36])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1701.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1702 (.D(key_mem_0__127__N_5088[37]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [37])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1702.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1703 (.D(key_mem_0__127__N_5088[38]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [38])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1703.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1704 (.D(key_mem_0__127__N_5088[39]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [39])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1704.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1705 (.D(key_mem_0__127__N_5088[40]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [40])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1705.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1706 (.D(key_mem_0__127__N_5088[41]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [41])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1706.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1707 (.D(key_mem_0__127__N_5088[42]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [42])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1707.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1708 (.D(key_mem_0__127__N_5088[43]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [43])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1708.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1709 (.D(key_mem_0__127__N_5088[44]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [44])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1709.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1710 (.D(key_mem_0__127__N_5088[45]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [45])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1710.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1711 (.D(key_mem_0__127__N_5088[46]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [46])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1711.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1712 (.D(key_mem_0__127__N_5088[47]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [47])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1712.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1713 (.D(key_mem_0__127__N_5088[48]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [48])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1713.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1714 (.D(key_mem_0__127__N_5088[49]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [49])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1714.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1715 (.D(key_mem_0__127__N_5088[50]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [50])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1715.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1716 (.D(key_mem_0__127__N_5088[51]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [51])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1716.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1717 (.D(key_mem_0__127__N_5088[52]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [52])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1717.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1718 (.D(key_mem_0__127__N_5088[53]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [53])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1718.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1719 (.D(key_mem_0__127__N_5088[54]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [54])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1719.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1720 (.D(key_mem_0__127__N_5088[55]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [55])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1720.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1721 (.D(key_mem_0__127__N_5088[56]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [56])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1721.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1722 (.D(key_mem_0__127__N_5088[57]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [57])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1722.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1723 (.D(key_mem_0__127__N_5088[58]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [58])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1723.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1724 (.D(key_mem_0__127__N_5088[59]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [59])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1724.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1725 (.D(key_mem_0__127__N_5088[60]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [60])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1725.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1726 (.D(key_mem_0__127__N_5088[61]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [61])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1726.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1727 (.D(key_mem_0__127__N_5088[62]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [62])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1727.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1728 (.D(key_mem_0__127__N_5088[63]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [63])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1728.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1729 (.D(key_mem_0__127__N_5088[64]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [64])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1729.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1730 (.D(key_mem_0__127__N_5088[65]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [65])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1730.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1731 (.D(key_mem_0__127__N_5088[66]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [66])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1731.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1732 (.D(key_mem_0__127__N_5088[67]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [67])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1732.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1733 (.D(key_mem_0__127__N_5088[68]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [68])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1733.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1734 (.D(key_mem_0__127__N_5088[69]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [69])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1734.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1735 (.D(key_mem_0__127__N_5088[70]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [70])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1735.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1736 (.D(key_mem_0__127__N_5088[71]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [71])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1736.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1737 (.D(key_mem_0__127__N_5088[72]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [72])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1737.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1738 (.D(key_mem_0__127__N_5088[73]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [73])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1738.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1739 (.D(key_mem_0__127__N_5088[74]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [74])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1739.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1740 (.D(key_mem_0__127__N_5088[75]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [75])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1740.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1741 (.D(key_mem_0__127__N_5088[76]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [76])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1741.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1742 (.D(key_mem_0__127__N_5088[77]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [77])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1742.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1743 (.D(key_mem_0__127__N_5088[78]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [78])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1743.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1744 (.D(key_mem_0__127__N_5088[79]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [79])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1744.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1745 (.D(key_mem_0__127__N_5088[80]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [80])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1745.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1746 (.D(key_mem_0__127__N_5088[81]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [81])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1746.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1747 (.D(key_mem_0__127__N_5088[82]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [82])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1747.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1748 (.D(key_mem_0__127__N_5088[83]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [83])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1748.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1749 (.D(key_mem_0__127__N_5088[84]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [84])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1749.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1750 (.D(key_mem_0__127__N_5088[85]), .SP(clk_c_enable_2136), 
            .CK(clk_c), .Q(\key_mem[1] [85])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1750.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1751 (.D(key_mem_0__127__N_5088[86]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[1] [86])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1751.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1752 (.D(key_mem_0__127__N_5088[87]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[1] [87])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1752.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1753 (.D(key_mem_0__127__N_5088[88]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[1] [88])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1753.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1754 (.D(key_mem_0__127__N_5088[89]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[1] [89])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1754.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1755 (.D(key_mem_0__127__N_5088[90]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[1] [90])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1755.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1756 (.D(key_mem_0__127__N_5088[91]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[1] [91])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1756.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1757 (.D(key_mem_0__127__N_5088[92]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[1] [92])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1757.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1758 (.D(key_mem_0__127__N_5088[93]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[1] [93])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1758.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1759 (.D(key_mem_0__127__N_5088[94]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[1] [94])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1759.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1760 (.D(key_mem_0__127__N_5088[95]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[1] [95])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1760.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1761 (.D(key_mem_0__127__N_5088[96]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[1] [96])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1761.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1762 (.D(key_mem_0__127__N_5088[97]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[1] [97])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1762.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1763 (.D(key_mem_0__127__N_5088[98]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[1] [98])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1763.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1764 (.D(key_mem_0__127__N_5088[99]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[1] [99])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1764.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1765 (.D(key_mem_0__127__N_5088[100]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[1] [100])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1765.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1766 (.D(key_mem_0__127__N_5088[101]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[1] [101])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1766.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1767 (.D(key_mem_0__127__N_5088[102]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[1] [102])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1767.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1768 (.D(key_mem_0__127__N_5088[103]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[1] [103])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1768.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1769 (.D(key_mem_0__127__N_5088[104]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[1] [104])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1769.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1770 (.D(key_mem_0__127__N_5088[105]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[1] [105])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1770.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1771 (.D(key_mem_0__127__N_5088[106]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[1] [106])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1771.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1772 (.D(key_mem_0__127__N_5088[107]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[1] [107])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1772.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1773 (.D(key_mem_0__127__N_5088[108]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[1] [108])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1773.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1774 (.D(key_mem_0__127__N_5088[109]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[1] [109])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1774.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1775 (.D(key_mem_0__127__N_5088[110]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[1] [110])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1775.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1776 (.D(key_mem_0__127__N_5088[111]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[1] [111])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1776.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1777 (.D(key_mem_0__127__N_5088[112]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[1] [112])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1777.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1778 (.D(key_mem_0__127__N_5088[113]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[1] [113])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1778.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1779 (.D(key_mem_0__127__N_5088[114]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[1] [114])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1779.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1780 (.D(key_mem_0__127__N_5088[115]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[1] [115])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1780.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1781 (.D(key_mem_0__127__N_5088[116]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[1] [116])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1781.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1782 (.D(key_mem_0__127__N_5088[117]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[1] [117])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1782.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1783 (.D(key_mem_0__127__N_5088[118]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[1] [118])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1783.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1784 (.D(key_mem_0__127__N_5088[119]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[1] [119])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1784.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1785 (.D(key_mem_0__127__N_5088[120]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[1] [120])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1785.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1786 (.D(key_mem_0__127__N_5088[121]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[1] [121])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1786.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1787 (.D(key_mem_0__127__N_5088[122]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[1] [122])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1787.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1788 (.D(key_mem_0__127__N_5088[123]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[1] [123])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1788.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1789 (.D(key_mem_0__127__N_5088[124]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[1] [124])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1789.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1790 (.D(key_mem_0__127__N_5088[125]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[1] [125])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1790.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1791 (.D(key_mem_0__127__N_5088[126]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[1] [126])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1791.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1792 (.D(key_mem_0__127__N_5088[127]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[1] [127])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1792.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1793 (.D(key_mem_0__127__N_4960[0]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[0] [0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1793.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1794 (.D(key_mem_0__127__N_4960[1]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[0] [1])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1794.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1795 (.D(key_mem_0__127__N_4960[2]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[0] [2])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1795.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1796 (.D(key_mem_0__127__N_4960[3]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[0] [3])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1796.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1797 (.D(key_mem_0__127__N_4960[4]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[0] [4])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1797.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1798 (.D(key_mem_0__127__N_4960[5]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[0] [5])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1798.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1799 (.D(key_mem_0__127__N_4960[6]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[0] [6])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1799.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1800 (.D(key_mem_0__127__N_4960[7]), .SP(clk_c_enable_2186), 
            .CK(clk_c), .Q(\key_mem[0] [7])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1800.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1801 (.D(key_mem_0__127__N_4960[8]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [8])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1801.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1802 (.D(key_mem_0__127__N_4960[9]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [9])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1802.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1803 (.D(key_mem_0__127__N_4960[10]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [10])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1803.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1804 (.D(key_mem_0__127__N_4960[11]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [11])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1804.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1805 (.D(key_mem_0__127__N_4960[12]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [12])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1805.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1806 (.D(key_mem_0__127__N_4960[13]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [13])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1806.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1807 (.D(key_mem_0__127__N_4960[14]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [14])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1807.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1808 (.D(key_mem_0__127__N_4960[15]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [15])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1808.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1809 (.D(key_mem_0__127__N_4960[16]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [16])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1809.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1810 (.D(key_mem_0__127__N_4960[17]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [17])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1810.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1811 (.D(key_mem_0__127__N_4960[18]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [18])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1811.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1812 (.D(key_mem_0__127__N_4960[19]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [19])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1812.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1813 (.D(key_mem_0__127__N_4960[20]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [20])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1813.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1814 (.D(key_mem_0__127__N_4960[21]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [21])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1814.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1815 (.D(key_mem_0__127__N_4960[22]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [22])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1815.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1816 (.D(key_mem_0__127__N_4960[23]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [23])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1816.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1817 (.D(key_mem_0__127__N_4960[24]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [24])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1817.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1818 (.D(key_mem_0__127__N_4960[25]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [25])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1818.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1819 (.D(key_mem_0__127__N_4960[26]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [26])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1819.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1820 (.D(key_mem_0__127__N_4960[27]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [27])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1820.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1821 (.D(key_mem_0__127__N_4960[28]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [28])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1821.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1822 (.D(key_mem_0__127__N_4960[29]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [29])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1822.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1823 (.D(key_mem_0__127__N_4960[30]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [30])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1823.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1824 (.D(key_mem_0__127__N_4960[31]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [31])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1824.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1825 (.D(key_mem_0__127__N_4960[32]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [32])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1825.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1826 (.D(key_mem_0__127__N_4960[33]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [33])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1826.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1827 (.D(key_mem_0__127__N_4960[34]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [34])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1827.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1828 (.D(key_mem_0__127__N_4960[35]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [35])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1828.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1829 (.D(key_mem_0__127__N_4960[36]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [36])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1829.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1830 (.D(key_mem_0__127__N_4960[37]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [37])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1830.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1831 (.D(key_mem_0__127__N_4960[38]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [38])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1831.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1832 (.D(key_mem_0__127__N_4960[39]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [39])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1832.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1833 (.D(key_mem_0__127__N_4960[40]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [40])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1833.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1834 (.D(key_mem_0__127__N_4960[41]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [41])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1834.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1835 (.D(key_mem_0__127__N_4960[42]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [42])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1835.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1836 (.D(key_mem_0__127__N_4960[43]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [43])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1836.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1837 (.D(key_mem_0__127__N_4960[44]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [44])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1837.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1838 (.D(key_mem_0__127__N_4960[45]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [45])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1838.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1839 (.D(key_mem_0__127__N_4960[46]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [46])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1839.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1840 (.D(key_mem_0__127__N_4960[47]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [47])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1840.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1841 (.D(key_mem_0__127__N_4960[48]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [48])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1841.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1842 (.D(key_mem_0__127__N_4960[49]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [49])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1842.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1843 (.D(key_mem_0__127__N_4960[50]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [50])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1843.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1844 (.D(key_mem_0__127__N_4960[51]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [51])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1844.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1845 (.D(key_mem_0__127__N_4960[52]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [52])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1845.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1846 (.D(key_mem_0__127__N_4960[53]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [53])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1846.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1847 (.D(key_mem_0__127__N_4960[54]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [54])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1847.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1848 (.D(key_mem_0__127__N_4960[55]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [55])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1848.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1849 (.D(key_mem_0__127__N_4960[56]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [56])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1849.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1850 (.D(key_mem_0__127__N_4960[57]), .SP(clk_c_enable_2236), 
            .CK(clk_c), .Q(\key_mem[0] [57])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1850.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1851 (.D(key_mem_0__127__N_4960[58]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [58])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1851.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1852 (.D(key_mem_0__127__N_4960[59]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [59])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1852.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1853 (.D(key_mem_0__127__N_4960[60]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [60])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1853.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1854 (.D(key_mem_0__127__N_4960[61]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [61])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1854.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1855 (.D(key_mem_0__127__N_4960[62]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [62])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1855.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1856 (.D(key_mem_0__127__N_4960[63]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [63])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1856.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1857 (.D(key_mem_0__127__N_4960[64]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [64])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1857.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1858 (.D(key_mem_0__127__N_4960[65]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [65])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1858.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1859 (.D(key_mem_0__127__N_4960[66]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [66])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1859.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1860 (.D(key_mem_0__127__N_4960[67]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [67])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1860.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1861 (.D(key_mem_0__127__N_4960[68]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [68])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1861.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1862 (.D(key_mem_0__127__N_4960[69]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [69])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1862.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1863 (.D(key_mem_0__127__N_4960[70]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [70])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1863.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1864 (.D(key_mem_0__127__N_4960[71]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [71])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1864.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1865 (.D(key_mem_0__127__N_4960[72]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [72])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1865.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1866 (.D(key_mem_0__127__N_4960[73]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [73])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1866.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1867 (.D(key_mem_0__127__N_4960[74]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [74])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1867.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1868 (.D(key_mem_0__127__N_4960[75]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [75])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1868.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1869 (.D(key_mem_0__127__N_4960[76]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [76])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1869.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1870 (.D(key_mem_0__127__N_4960[77]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [77])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1870.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1871 (.D(key_mem_0__127__N_4960[78]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [78])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1871.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1872 (.D(key_mem_0__127__N_4960[79]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [79])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1872.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1873 (.D(key_mem_0__127__N_4960[80]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [80])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1873.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1874 (.D(key_mem_0__127__N_4960[81]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [81])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1874.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1875 (.D(key_mem_0__127__N_4960[82]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [82])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1875.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1876 (.D(key_mem_0__127__N_4960[83]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [83])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1876.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1877 (.D(key_mem_0__127__N_4960[84]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [84])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1877.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1878 (.D(key_mem_0__127__N_4960[85]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [85])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1878.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1879 (.D(key_mem_0__127__N_4960[86]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [86])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1879.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1880 (.D(key_mem_0__127__N_4960[87]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [87])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1880.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1881 (.D(key_mem_0__127__N_4960[88]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [88])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1881.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1882 (.D(key_mem_0__127__N_4960[89]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [89])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1882.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1883 (.D(key_mem_0__127__N_4960[90]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [90])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1883.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1884 (.D(key_mem_0__127__N_4960[91]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [91])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1884.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1885 (.D(key_mem_0__127__N_4960[92]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [92])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1885.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1886 (.D(key_mem_0__127__N_4960[93]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [93])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1886.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1887 (.D(key_mem_0__127__N_4960[94]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [94])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1887.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1888 (.D(key_mem_0__127__N_4960[95]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [95])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1888.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1889 (.D(key_mem_0__127__N_4960[96]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [96])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1889.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1890 (.D(key_mem_0__127__N_4960[97]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [97])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1890.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1891 (.D(key_mem_0__127__N_4960[98]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [98])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1891.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1892 (.D(key_mem_0__127__N_4960[99]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [99])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1892.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1893 (.D(key_mem_0__127__N_4960[100]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [100])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1893.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1894 (.D(key_mem_0__127__N_4960[101]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [101])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1894.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1895 (.D(key_mem_0__127__N_4960[102]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [102])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1895.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1896 (.D(key_mem_0__127__N_4960[103]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [103])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1896.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1897 (.D(key_mem_0__127__N_4960[104]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [104])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1897.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1898 (.D(key_mem_0__127__N_4960[105]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [105])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1898.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1899 (.D(key_mem_0__127__N_4960[106]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [106])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1899.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1900 (.D(key_mem_0__127__N_4960[107]), .SP(clk_c_enable_2286), 
            .CK(clk_c), .Q(\key_mem[0] [107])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1900.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1901 (.D(key_mem_0__127__N_4960[108]), .SP(n6361[1]), 
            .CK(clk_c), .Q(\key_mem[0] [108])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1901.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1902 (.D(key_mem_0__127__N_4960[109]), .SP(n6361[1]), 
            .CK(clk_c), .Q(\key_mem[0] [109])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1902.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1903 (.D(key_mem_0__127__N_4960[110]), .SP(n6361[1]), 
            .CK(clk_c), .Q(\key_mem[0] [110])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1903.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1904 (.D(key_mem_0__127__N_4960[111]), .SP(n6361[1]), 
            .CK(clk_c), .Q(\key_mem[0] [111])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1904.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1905 (.D(key_mem_0__127__N_4960[112]), .SP(n6361[1]), 
            .CK(clk_c), .Q(\key_mem[0] [112])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1905.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1906 (.D(key_mem_0__127__N_4960[113]), .SP(n6361[1]), 
            .CK(clk_c), .Q(\key_mem[0] [113])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1906.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1907 (.D(key_mem_0__127__N_4960[114]), .SP(n6361[1]), 
            .CK(clk_c), .Q(\key_mem[0] [114])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1907.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1908 (.D(key_mem_0__127__N_4960[115]), .SP(n6361[1]), 
            .CK(clk_c), .Q(\key_mem[0] [115])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1908.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1909 (.D(key_mem_0__127__N_4960[116]), .SP(n6361[1]), 
            .CK(clk_c), .Q(\key_mem[0] [116])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1909.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1910 (.D(key_mem_0__127__N_4960[117]), .SP(n6361[1]), 
            .CK(clk_c), .Q(\key_mem[0] [117])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1910.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1911 (.D(key_mem_0__127__N_4960[118]), .SP(n6361[1]), 
            .CK(clk_c), .Q(\key_mem[0] [118])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1911.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1912 (.D(key_mem_0__127__N_4960[119]), .SP(n6361[1]), 
            .CK(clk_c), .Q(\key_mem[0] [119])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1912.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1913 (.D(key_mem_0__127__N_4960[120]), .SP(n6361[1]), 
            .CK(clk_c), .Q(\key_mem[0] [120])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1913.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1914 (.D(key_mem_0__127__N_4960[121]), .SP(n6361[1]), 
            .CK(clk_c), .Q(\key_mem[0] [121])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1914.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1915 (.D(key_mem_0__127__N_4960[122]), .SP(n6361[1]), 
            .CK(clk_c), .Q(\key_mem[0] [122])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1915.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1916 (.D(key_mem_0__127__N_4960[123]), .SP(n6361[1]), 
            .CK(clk_c), .Q(\key_mem[0] [123])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1916.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1917 (.D(key_mem_0__127__N_4960[124]), .SP(n6361[1]), 
            .CK(clk_c), .Q(\key_mem[0] [124])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1917.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1918 (.D(key_mem_0__127__N_4960[125]), .SP(n6361[1]), 
            .CK(clk_c), .Q(\key_mem[0] [125])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1918.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1919 (.D(key_mem_0__127__N_4960[126]), .SP(n6361[1]), 
            .CK(clk_c), .Q(\key_mem[0] [126])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1919.GSR = "ENABLED";
    FD1P3AX key_mem_14___i1920 (.D(key_mem_0__127__N_4960[127]), .SP(n6361[1]), 
            .CK(clk_c), .Q(\key_mem[0] [127])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam key_mem_14___i1920.GSR = "ENABLED";
    FD1P3IX prev_key1_reg__i2 (.D(\prev_key1_new_127__N_4787[1] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(keymem_sboxw[1])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i2.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i3 (.D(\prev_key1_new_127__N_4787[2] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(keymem_sboxw[2])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i3.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i4 (.D(\prev_key1_new_127__N_4787[3] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(keymem_sboxw[3])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i4.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i5 (.D(\prev_key1_new_127__N_4787[4] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(keymem_sboxw[4])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i5.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i6 (.D(\prev_key1_new_127__N_4787[5] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(keymem_sboxw[5])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i6.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i7 (.D(\prev_key1_new_127__N_4787[6] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(keymem_sboxw[6])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i7.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i8 (.D(\prev_key1_new_127__N_4787[7] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(keymem_sboxw[7])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i8.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i9 (.D(\prev_key1_new_127__N_4787[8] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(keymem_sboxw[8])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i9.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i10 (.D(\prev_key1_new_127__N_4787[9] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(keymem_sboxw[9])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i10.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i11 (.D(\prev_key1_new_127__N_4787[10] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(keymem_sboxw[10])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i11.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i12 (.D(\prev_key1_new_127__N_4787[11] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(keymem_sboxw[11])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i12.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i13 (.D(\prev_key1_new_127__N_4787[12] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(keymem_sboxw[12])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i13.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i14 (.D(\prev_key1_new_127__N_4787[13] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(keymem_sboxw[13])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i14.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i15 (.D(\prev_key1_new_127__N_4787[14] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(keymem_sboxw[14])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i15.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i16 (.D(\prev_key1_new_127__N_4787[15] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(keymem_sboxw[15])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i16.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i17 (.D(\prev_key1_new_127__N_4787[16] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(keymem_sboxw[16])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i17.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i18 (.D(\prev_key1_new_127__N_4787[17] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(keymem_sboxw[17])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i18.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i19 (.D(\prev_key1_new_127__N_4787[18] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(keymem_sboxw[18])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i19.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i20 (.D(\prev_key1_new_127__N_4787[19] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(keymem_sboxw[19])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i20.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i21 (.D(\prev_key1_new_127__N_4787[20] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(keymem_sboxw[20])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i21.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i22 (.D(\prev_key1_new_127__N_4787[21] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(keymem_sboxw[21])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i22.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i23 (.D(\prev_key1_new_127__N_4787[22] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(keymem_sboxw[22])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i23.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i24 (.D(\prev_key1_new_127__N_4787[23] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(keymem_sboxw[23])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i24.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i25 (.D(\prev_key1_new_127__N_4787[24] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(keymem_sboxw[24])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i25.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i26 (.D(\prev_key1_new_127__N_4787[25] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(keymem_sboxw[25])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i26.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i27 (.D(\prev_key1_new_127__N_4787[26] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(keymem_sboxw[26])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i27.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i28 (.D(\prev_key1_new_127__N_4787[27] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(keymem_sboxw[27])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i28.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i29 (.D(\prev_key1_new_127__N_4787[28] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(keymem_sboxw[28])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i29.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i30 (.D(\prev_key1_new_127__N_4787[29] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(keymem_sboxw[29])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i30.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i31 (.D(\prev_key1_new_127__N_4787[30] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(keymem_sboxw[30])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i31.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i32 (.D(\prev_key1_new_127__N_4787[31] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(keymem_sboxw[31])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i32.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i33 (.D(\prev_key1_new_127__N_4787[32] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[32])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i33.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i34 (.D(\prev_key1_new_127__N_4787[33] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[33])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i34.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i35 (.D(\prev_key1_new_127__N_4787[34] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[34])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i35.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i36 (.D(\prev_key1_new_127__N_4787[35] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[35])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i36.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i37 (.D(\prev_key1_new_127__N_4787[36] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[36])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i37.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i38 (.D(\prev_key1_new_127__N_4787[37] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[37])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i38.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i39 (.D(\prev_key1_new_127__N_4787[38] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[38])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i39.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i40 (.D(\prev_key1_new_127__N_4787[39] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[39])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i40.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i41 (.D(\prev_key1_new_127__N_4787[40] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[40])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i41.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i42 (.D(\prev_key1_new_127__N_4787[41] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[41])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i42.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i43 (.D(\prev_key1_new_127__N_4787[42] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[42])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i43.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i44 (.D(\prev_key1_new_127__N_4787[43] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[43])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i44.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i45 (.D(\prev_key1_new_127__N_4787[44] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[44])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i45.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i46 (.D(\prev_key1_new_127__N_4787[45] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[45])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i46.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i47 (.D(\prev_key1_new_127__N_4787[46] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[46])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i47.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i48 (.D(\prev_key1_new_127__N_4787[47] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[47])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i48.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i49 (.D(\prev_key1_new_127__N_4787[48] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[48])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i49.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i50 (.D(\prev_key1_new_127__N_4787[49] ), .SP(clk_c_enable_2335), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[49])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i50.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i51 (.D(\prev_key1_new_127__N_4787[50] ), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[50])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i51.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i52 (.D(\prev_key1_new_127__N_4787[51] ), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[51])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i52.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i53 (.D(\prev_key1_new_127__N_4787[52] ), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[52])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i53.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i54 (.D(\prev_key1_new_127__N_4787[53] ), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[53])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i54.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i55 (.D(\prev_key1_new_127__N_4787[54] ), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[54])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i55.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i56 (.D(\prev_key1_new_127__N_4787[55] ), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[55])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i56.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i57 (.D(\prev_key1_new_127__N_4787[56] ), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[56])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i57.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i58 (.D(\prev_key1_new_127__N_4787[57] ), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[57])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i58.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i59 (.D(\prev_key1_new_127__N_4787[58] ), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[58])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i59.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i60 (.D(\prev_key1_new_127__N_4787[59] ), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[59])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i60.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i61 (.D(\prev_key1_new_127__N_4787[60] ), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[60])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i61.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i62 (.D(\prev_key1_new_127__N_4787[61] ), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[61])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i62.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i63 (.D(\prev_key1_new_127__N_4787[62] ), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[62])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i63.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i64 (.D(\prev_key1_new_127__N_4787[63] ), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[63])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i64.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i65 (.D(prev_key1_new_127__N_4787[64]), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[64])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i65.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i66 (.D(prev_key1_new_127__N_4787[65]), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[65])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i66.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i67 (.D(prev_key1_new_127__N_4787[66]), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[66])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i67.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i68 (.D(prev_key1_new_127__N_4787[67]), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[67])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i68.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i69 (.D(prev_key1_new_127__N_4787[68]), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[68])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i69.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i70 (.D(prev_key1_new_127__N_4787[69]), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[69])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i70.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i71 (.D(prev_key1_new_127__N_4787[70]), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[70])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i71.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i72 (.D(prev_key1_new_127__N_4787[71]), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[71])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i72.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i73 (.D(prev_key1_new_127__N_4787[72]), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[72])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i73.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i74 (.D(prev_key1_new_127__N_4787[73]), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[73])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i74.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i75 (.D(prev_key1_new_127__N_4787[74]), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[74])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i75.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i76 (.D(prev_key1_new_127__N_4787[75]), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[75])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i76.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i77 (.D(prev_key1_new_127__N_4787[76]), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[76])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i77.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i78 (.D(prev_key1_new_127__N_4787[77]), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[77])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i78.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i79 (.D(prev_key1_new_127__N_4787[78]), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[78])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i79.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i80 (.D(prev_key1_new_127__N_4787[79]), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[79])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i80.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i81 (.D(prev_key1_new_127__N_4787[80]), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[80])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i81.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i82 (.D(prev_key1_new_127__N_4787[81]), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[81])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i82.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i83 (.D(prev_key1_new_127__N_4787[82]), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[82])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i83.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i84 (.D(prev_key1_new_127__N_4787[83]), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[83])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i84.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i85 (.D(prev_key1_new_127__N_4787[84]), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[84])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i85.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i86 (.D(prev_key1_new_127__N_4787[85]), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[85])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i86.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i87 (.D(prev_key1_new_127__N_4787[86]), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[86])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i87.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i88 (.D(prev_key1_new_127__N_4787[87]), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[87])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i88.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i89 (.D(prev_key1_new_127__N_4787[88]), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[88])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i89.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i90 (.D(prev_key1_new_127__N_4787[89]), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[89])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i90.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i91 (.D(prev_key1_new_127__N_4787[90]), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[90])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i91.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i92 (.D(prev_key1_new_127__N_4787[91]), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[91])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i92.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i93 (.D(prev_key1_new_127__N_4787[92]), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[92])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i93.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i94 (.D(prev_key1_new_127__N_4787[93]), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[93])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i94.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i95 (.D(prev_key1_new_127__N_4787[94]), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[94])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i95.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i96 (.D(prev_key1_new_127__N_4787[95]), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[95])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i96.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i97 (.D(prev_key1_new_127__N_4787[96]), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[96])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i97.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i98 (.D(prev_key1_new_127__N_4787[97]), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[97])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i98.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i99 (.D(prev_key1_new_127__N_4787[98]), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[98])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i99.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i100 (.D(prev_key1_new_127__N_4787[99]), .SP(clk_c_enable_2385), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[99])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i100.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i101 (.D(prev_key1_new_127__N_4787[100]), .SP(clk_c_enable_2413), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[100])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i101.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i102 (.D(prev_key1_new_127__N_4787[101]), .SP(clk_c_enable_2413), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[101])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i102.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i103 (.D(prev_key1_new_127__N_4787[102]), .SP(clk_c_enable_2413), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[102])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i103.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i104 (.D(prev_key1_new_127__N_4787[103]), .SP(clk_c_enable_2413), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[103])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i104.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i105 (.D(prev_key1_new_127__N_4787[104]), .SP(clk_c_enable_2413), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[104])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i105.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i106 (.D(prev_key1_new_127__N_4787[105]), .SP(clk_c_enable_2413), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[105])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i106.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i107 (.D(prev_key1_new_127__N_4787[106]), .SP(clk_c_enable_2413), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[106])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i107.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i108 (.D(prev_key1_new_127__N_4787[107]), .SP(clk_c_enable_2413), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[107])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i108.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i109 (.D(prev_key1_new_127__N_4787[108]), .SP(clk_c_enable_2413), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[108])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i109.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i110 (.D(prev_key1_new_127__N_4787[109]), .SP(clk_c_enable_2413), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[109])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i110.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i111 (.D(prev_key1_new_127__N_4787[110]), .SP(clk_c_enable_2413), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[110])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i111.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i112 (.D(prev_key1_new_127__N_4787[111]), .SP(clk_c_enable_2413), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[111])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i112.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i113 (.D(prev_key1_new_127__N_4787[112]), .SP(clk_c_enable_2413), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[112])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i113.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i114 (.D(prev_key1_new_127__N_4787[113]), .SP(clk_c_enable_2413), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[113])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i114.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i115 (.D(prev_key1_new_127__N_4787[114]), .SP(clk_c_enable_2413), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[114])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i115.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i116 (.D(prev_key1_new_127__N_4787[115]), .SP(clk_c_enable_2413), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[115])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i116.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i117 (.D(prev_key1_new_127__N_4787[116]), .SP(clk_c_enable_2413), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[116])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i117.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i118 (.D(prev_key1_new_127__N_4787[117]), .SP(clk_c_enable_2413), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[117])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i118.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i119 (.D(prev_key1_new_127__N_4787[118]), .SP(clk_c_enable_2413), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[118])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i119.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i120 (.D(prev_key1_new_127__N_4787[119]), .SP(clk_c_enable_2413), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[119])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i120.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i121 (.D(prev_key1_new_127__N_4787[120]), .SP(clk_c_enable_2413), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[120])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i121.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i122 (.D(prev_key1_new_127__N_4787[121]), .SP(clk_c_enable_2413), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[121])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i122.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i123 (.D(prev_key1_new_127__N_4787[122]), .SP(clk_c_enable_2413), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[122])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i123.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i124 (.D(prev_key1_new_127__N_4787[123]), .SP(clk_c_enable_2413), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[123])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i124.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i125 (.D(prev_key1_new_127__N_4787[124]), .SP(clk_c_enable_2413), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[124])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i125.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i126 (.D(prev_key1_new_127__N_4787[125]), .SP(clk_c_enable_2413), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[125])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i126.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i127 (.D(prev_key1_new_127__N_4787[126]), .SP(clk_c_enable_2413), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[126])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i127.GSR = "DISABLED";
    FD1P3IX prev_key1_reg__i128 (.D(prev_key1_new_127__N_4787[127]), .SP(clk_c_enable_2413), 
            .CD(GND_net), .CK(clk_c), .Q(prev_key1_reg[127])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam prev_key1_reg__i128.GSR = "DISABLED";
    LUT4 mux_20_i3_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [2]), 
         .D(key_mem_new[2]), .Z(key_mem_0__127__N_5344[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i3_3_lut_4_lut.init = 16'hf2d0;
    L6MUX21 i25441 (.D0(n30597), .D1(n33431), .SD(\muxed_round_nr[2] ), 
            .Z(n30600));
    L6MUX21 i25447 (.D0(n30602), .D1(n30603), .SD(\muxed_round_nr[2] ), 
            .Z(n30606));
    L6MUX21 i25448 (.D0(n30604), .D1(n33432), .SD(\muxed_round_nr[2] ), 
            .Z(n30607));
    LUT4 round_3__I_0_Mux_103_i11_3_lut (.A(\key_mem[12] [103]), .B(\key_mem[13] [103]), 
         .C(n33952), .Z(n11_adj_123)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_103_i11_3_lut.init = 16'hcaca;
    L6MUX21 i25454 (.D0(n30609), .D1(n30610), .SD(\muxed_round_nr[2] ), 
            .Z(n30613));
    LUT4 mux_20_i4_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [3]), 
         .D(key_mem_new[3]), .Z(key_mem_0__127__N_5344[3])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i4_3_lut_4_lut.init = 16'hf2d0;
    L6MUX21 i25455 (.D0(n30611), .D1(n33433), .SD(\muxed_round_nr[2] ), 
            .Z(n30614));
    LUT4 mux_20_i5_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [4]), 
         .D(key_mem_new[4]), .Z(key_mem_0__127__N_5344[4])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i5_3_lut_4_lut.init = 16'hf2d0;
    L6MUX21 i25461 (.D0(n30616), .D1(n30617), .SD(\muxed_round_nr[2] ), 
            .Z(n30620));
    LUT4 mux_20_i6_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [5]), 
         .D(key_mem_new[5]), .Z(key_mem_0__127__N_5344[5])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i6_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i7_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [6]), 
         .D(key_mem_new[6]), .Z(key_mem_0__127__N_5344[6])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i7_3_lut_4_lut.init = 16'hf2d0;
    L6MUX21 i25462 (.D0(n30618), .D1(n33434), .SD(\muxed_round_nr[2] ), 
            .Z(n30621));
    LUT4 mux_20_i8_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [7]), 
         .D(key_mem_new[7]), .Z(key_mem_0__127__N_5344[7])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i8_3_lut_4_lut.init = 16'hf2d0;
    LUT4 round_3__I_0_Mux_103_i9_3_lut (.A(\key_mem[10] [103]), .B(\key_mem[11] [103]), 
         .C(n33952), .Z(n9_adj_9254)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_103_i9_3_lut.init = 16'hcaca;
    LUT4 mux_20_i9_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [8]), 
         .D(key_mem_new[8]), .Z(key_mem_0__127__N_5344[8])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i9_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i10_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [9]), 
         .D(key_mem_new[9]), .Z(key_mem_0__127__N_5344[9])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i10_3_lut_4_lut.init = 16'hf2d0;
    LUT4 round_3__I_0_Mux_103_i8_3_lut (.A(\key_mem[8] [103]), .B(\key_mem[9] [103]), 
         .C(n33952), .Z(n8_adj_9255)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_103_i8_3_lut.init = 16'hcaca;
    L6MUX21 i25468 (.D0(n30623), .D1(n30624), .SD(\muxed_round_nr[2] ), 
            .Z(n30627));
    LUT4 mux_20_i11_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [10]), 
         .D(key_mem_new[10]), .Z(key_mem_0__127__N_5344[10])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i11_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i12_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [11]), 
         .D(key_mem_new[11]), .Z(key_mem_0__127__N_5344[11])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i12_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i13_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [12]), 
         .D(key_mem_new[12]), .Z(key_mem_0__127__N_5344[12])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i13_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i14_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [13]), 
         .D(key_mem_new[13]), .Z(key_mem_0__127__N_5344[13])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i14_3_lut_4_lut.init = 16'hf2d0;
    L6MUX21 i25469 (.D0(n30625), .D1(n33436), .SD(\muxed_round_nr[2] ), 
            .Z(n30628));
    L6MUX21 i25475 (.D0(n30630), .D1(n30631), .SD(\muxed_round_nr[2] ), 
            .Z(n30634));
    LUT4 mux_20_i15_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [14]), 
         .D(key_mem_new[14]), .Z(key_mem_0__127__N_5344[14])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i15_3_lut_4_lut.init = 16'hf2d0;
    L6MUX21 i25476 (.D0(n30632), .D1(n33441), .SD(\muxed_round_nr[2] ), 
            .Z(n30635));
    LUT4 mux_20_i16_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [15]), 
         .D(key_mem_new[15]), .Z(key_mem_0__127__N_5344[15])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i16_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i17_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [16]), 
         .D(key_mem_new[16]), .Z(key_mem_0__127__N_5344[16])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i17_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i18_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [17]), 
         .D(key_mem_new[17]), .Z(key_mem_0__127__N_5344[17])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i18_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i19_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [18]), 
         .D(key_mem_new[18]), .Z(key_mem_0__127__N_5344[18])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i19_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i20_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [19]), 
         .D(key_mem_new[19]), .Z(key_mem_0__127__N_5344[19])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i20_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i21_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [20]), 
         .D(key_mem_new[20]), .Z(key_mem_0__127__N_5344[20])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i21_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i22_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [21]), 
         .D(key_mem_new[21]), .Z(key_mem_0__127__N_5344[21])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i22_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i23_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [22]), 
         .D(key_mem_new[22]), .Z(key_mem_0__127__N_5344[22])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i23_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i24_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [23]), 
         .D(key_mem_new[23]), .Z(key_mem_0__127__N_5344[23])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i24_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i25_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [24]), 
         .D(key_mem_new[24]), .Z(key_mem_0__127__N_5344[24])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i25_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i26_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [25]), 
         .D(key_mem_new[25]), .Z(key_mem_0__127__N_5344[25])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i26_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i27_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [26]), 
         .D(key_mem_new[26]), .Z(key_mem_0__127__N_5344[26])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i27_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i28_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [27]), 
         .D(key_mem_new[27]), .Z(key_mem_0__127__N_5344[27])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i28_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i29_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [28]), 
         .D(key_mem_new[28]), .Z(key_mem_0__127__N_5344[28])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i29_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i30_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [29]), 
         .D(key_mem_new[29]), .Z(key_mem_0__127__N_5344[29])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i30_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i31_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [30]), 
         .D(key_mem_new[30]), .Z(key_mem_0__127__N_5344[30])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i31_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i32_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [31]), 
         .D(key_mem_new[31]), .Z(key_mem_0__127__N_5344[31])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i32_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i33_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [32]), 
         .D(key_mem_new[32]), .Z(key_mem_0__127__N_5344[32])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i33_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i34_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [33]), 
         .D(key_mem_new[33]), .Z(key_mem_0__127__N_5344[33])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i34_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i35_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [34]), 
         .D(key_mem_new[34]), .Z(key_mem_0__127__N_5344[34])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i35_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i36_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [35]), 
         .D(key_mem_new[35]), .Z(key_mem_0__127__N_5344[35])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i36_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i37_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [36]), 
         .D(key_mem_new[36]), .Z(key_mem_0__127__N_5344[36])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i37_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i38_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [37]), 
         .D(key_mem_new[37]), .Z(key_mem_0__127__N_5344[37])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i38_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i39_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [38]), 
         .D(key_mem_new[38]), .Z(key_mem_0__127__N_5344[38])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i39_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i40_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [39]), 
         .D(key_mem_new[39]), .Z(key_mem_0__127__N_5344[39])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i40_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i41_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [40]), 
         .D(key_mem_new[40]), .Z(key_mem_0__127__N_5344[40])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i41_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i42_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [41]), 
         .D(key_mem_new[41]), .Z(key_mem_0__127__N_5344[41])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i42_3_lut_4_lut.init = 16'hf2d0;
    LUT4 round_3__I_0_Mux_116_i5_3_lut (.A(\key_mem[6] [116]), .B(\key_mem[7] [116]), 
         .C(n33952), .Z(n5_adj_8957)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_116_i5_3_lut.init = 16'hcaca;
    LUT4 mux_20_i43_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [42]), 
         .D(key_mem_new[42]), .Z(key_mem_0__127__N_5344[42])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i43_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i44_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [43]), 
         .D(key_mem_new[43]), .Z(key_mem_0__127__N_5344[43])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i44_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i45_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [44]), 
         .D(key_mem_new[44]), .Z(key_mem_0__127__N_5344[44])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i45_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i46_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [45]), 
         .D(key_mem_new[45]), .Z(key_mem_0__127__N_5344[45])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i46_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i47_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [46]), 
         .D(key_mem_new[46]), .Z(key_mem_0__127__N_5344[46])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i47_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i48_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [47]), 
         .D(key_mem_new[47]), .Z(key_mem_0__127__N_5344[47])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i48_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i49_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [48]), 
         .D(key_mem_new[48]), .Z(key_mem_0__127__N_5344[48])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i49_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i50_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [49]), 
         .D(key_mem_new[49]), .Z(key_mem_0__127__N_5344[49])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i50_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i51_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [50]), 
         .D(key_mem_new[50]), .Z(key_mem_0__127__N_5344[50])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i51_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i52_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [51]), 
         .D(key_mem_new[51]), .Z(key_mem_0__127__N_5344[51])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i52_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i53_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [52]), 
         .D(key_mem_new[52]), .Z(key_mem_0__127__N_5344[52])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i53_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i54_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [53]), 
         .D(key_mem_new[53]), .Z(key_mem_0__127__N_5344[53])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i54_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i55_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [54]), 
         .D(key_mem_new[54]), .Z(key_mem_0__127__N_5344[54])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i55_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i56_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [55]), 
         .D(key_mem_new[55]), .Z(key_mem_0__127__N_5344[55])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i56_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i57_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [56]), 
         .D(key_mem_new[56]), .Z(key_mem_0__127__N_5344[56])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i57_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i58_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [57]), 
         .D(key_mem_new[57]), .Z(key_mem_0__127__N_5344[57])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i58_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i11_4_lut_adj_654 (.A(n5), .B(keymem_sboxw[24]), .C(init_state), 
         .D(n10_adj_9256), .Z(muxed_sboxw[24])) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(181[17:28])
    defparam i11_4_lut_adj_654.init = 16'hc5c0;
    LUT4 mux_20_i59_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [58]), 
         .D(key_mem_new[58]), .Z(key_mem_0__127__N_5344[58])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i59_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i60_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [59]), 
         .D(key_mem_new[59]), .Z(key_mem_0__127__N_5344[59])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i60_3_lut_4_lut.init = 16'hf2d0;
    L6MUX21 i25482 (.D0(n30637), .D1(n30638), .SD(\muxed_round_nr[2] ), 
            .Z(n30641));
    LUT4 mux_20_i61_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [60]), 
         .D(key_mem_new[60]), .Z(key_mem_0__127__N_5344[60])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i61_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i62_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [61]), 
         .D(key_mem_new[61]), .Z(key_mem_0__127__N_5344[61])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i62_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i63_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [62]), 
         .D(key_mem_new[62]), .Z(key_mem_0__127__N_5344[62])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i63_3_lut_4_lut.init = 16'hf2d0;
    LUT4 round_3__I_0_Mux_103_i5_3_lut (.A(\key_mem[6] [103]), .B(\key_mem[7] [103]), 
         .C(n33952), .Z(n5_adj_9257)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_103_i5_3_lut.init = 16'hcaca;
    L6MUX21 i25483 (.D0(n30639), .D1(n33446), .SD(\muxed_round_nr[2] ), 
            .Z(n30642));
    L6MUX21 i25489 (.D0(n30644), .D1(n30645), .SD(\muxed_round_nr[2] ), 
            .Z(n30648));
    L6MUX21 i25490 (.D0(n30646), .D1(n33448), .SD(\muxed_round_nr[2] ), 
            .Z(n30649));
    LUT4 mux_20_i64_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [63]), 
         .D(key_mem_new[63]), .Z(key_mem_0__127__N_5344[63])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i64_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i11_4_lut_adj_655 (.A(n5), .B(keymem_sboxw[25]), .C(init_state), 
         .D(n10_adj_9258), .Z(muxed_sboxw[25])) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(181[17:28])
    defparam i11_4_lut_adj_655.init = 16'hc5c0;
    LUT4 mux_20_i65_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [64]), 
         .D(key_mem_new[64]), .Z(key_mem_0__127__N_5344[64])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i65_3_lut_4_lut.init = 16'hf2d0;
    LUT4 round_3__I_0_Mux_103_i4_3_lut (.A(\key_mem[4] [103]), .B(\key_mem[5] [103]), 
         .C(n33952), .Z(n4_adj_9259)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_103_i4_3_lut.init = 16'hcaca;
    LUT4 mux_20_i66_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [65]), 
         .D(key_mem_new[65]), .Z(key_mem_0__127__N_5344[65])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i66_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i67_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [66]), 
         .D(key_mem_new[66]), .Z(key_mem_0__127__N_5344[66])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i67_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i68_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [67]), 
         .D(key_mem_new[67]), .Z(key_mem_0__127__N_5344[67])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i68_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i69_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [68]), 
         .D(key_mem_new[68]), .Z(key_mem_0__127__N_5344[68])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i69_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i70_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [69]), 
         .D(key_mem_new[69]), .Z(key_mem_0__127__N_5344[69])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i70_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i71_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [70]), 
         .D(key_mem_new[70]), .Z(key_mem_0__127__N_5344[70])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i71_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i72_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [71]), 
         .D(key_mem_new[71]), .Z(key_mem_0__127__N_5344[71])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i72_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i73_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [72]), 
         .D(key_mem_new[72]), .Z(key_mem_0__127__N_5344[72])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i73_3_lut_4_lut.init = 16'hf2d0;
    L6MUX21 i25496 (.D0(n30651), .D1(n30652), .SD(\muxed_round_nr[2] ), 
            .Z(n30655));
    LUT4 mux_20_i74_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [73]), 
         .D(key_mem_new[73]), .Z(key_mem_0__127__N_5344[73])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i74_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i75_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [74]), 
         .D(key_mem_new[74]), .Z(key_mem_0__127__N_5344[74])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i75_3_lut_4_lut.init = 16'hf2d0;
    L6MUX21 i25497 (.D0(n30653), .D1(n33449), .SD(\muxed_round_nr[2] ), 
            .Z(n30656));
    LUT4 mux_20_i76_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [75]), 
         .D(key_mem_new[75]), .Z(key_mem_0__127__N_5344[75])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i76_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i77_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [76]), 
         .D(key_mem_new[76]), .Z(key_mem_0__127__N_5344[76])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i77_3_lut_4_lut.init = 16'hf2d0;
    L6MUX21 i25503 (.D0(n30658), .D1(n30659), .SD(\muxed_round_nr[2] ), 
            .Z(n30662));
    LUT4 mux_20_i78_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [77]), 
         .D(key_mem_new[77]), .Z(key_mem_0__127__N_5344[77])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i78_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i11_4_lut_adj_656 (.A(n5), .B(keymem_sboxw[26]), .C(init_state), 
         .D(n10_adj_9260), .Z(muxed_sboxw[26])) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(181[17:28])
    defparam i11_4_lut_adj_656.init = 16'hc5c0;
    L6MUX21 i25504 (.D0(n30660), .D1(n33450), .SD(\muxed_round_nr[2] ), 
            .Z(n30663));
    LUT4 mux_20_i79_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [78]), 
         .D(key_mem_new[78]), .Z(key_mem_0__127__N_5344[78])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i79_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i11_4_lut_adj_657 (.A(n5), .B(keymem_sboxw[27]), .C(init_state), 
         .D(n10_adj_9261), .Z(muxed_sboxw[27])) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(181[17:28])
    defparam i11_4_lut_adj_657.init = 16'hc5c0;
    L6MUX21 i25510 (.D0(n30665), .D1(n30666), .SD(\muxed_round_nr[2] ), 
            .Z(n30669));
    LUT4 mux_20_i80_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [79]), 
         .D(key_mem_new[79]), .Z(key_mem_0__127__N_5344[79])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i80_3_lut_4_lut.init = 16'hf2d0;
    L6MUX21 i25511 (.D0(n30667), .D1(n33451), .SD(\muxed_round_nr[2] ), 
            .Z(n30670));
    LUT4 mux_20_i81_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [80]), 
         .D(key_mem_new[80]), .Z(key_mem_0__127__N_5344[80])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i81_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i82_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [81]), 
         .D(key_mem_new[81]), .Z(key_mem_0__127__N_5344[81])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i82_3_lut_4_lut.init = 16'hf2d0;
    LUT4 round_3__I_0_Mux_103_i2_3_lut (.A(\key_mem[2] [103]), .B(\key_mem[3] [103]), 
         .C(n33952), .Z(n2_adj_9262)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_103_i2_3_lut.init = 16'hcaca;
    L6MUX21 i25517 (.D0(n30672), .D1(n30673), .SD(\muxed_round_nr[2] ), 
            .Z(n30676));
    LUT4 mux_20_i83_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [82]), 
         .D(key_mem_new[82]), .Z(key_mem_0__127__N_5344[82])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i83_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i84_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [83]), 
         .D(key_mem_new[83]), .Z(key_mem_0__127__N_5344[83])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i84_3_lut_4_lut.init = 16'hf2d0;
    LUT4 round_3__I_0_Mux_103_i1_3_lut (.A(\key_mem[0] [103]), .B(\key_mem[1] [103]), 
         .C(n33952), .Z(n1_adj_9263)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_103_i1_3_lut.init = 16'hcaca;
    L6MUX21 i25518 (.D0(n30674), .D1(n33452), .SD(\muxed_round_nr[2] ), 
            .Z(n30677));
    LUT4 mux_20_i85_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [84]), 
         .D(key_mem_new[84]), .Z(key_mem_0__127__N_5344[84])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i85_3_lut_4_lut.init = 16'hf2d0;
    L6MUX21 i25524 (.D0(n30679), .D1(n30680), .SD(\muxed_round_nr[2] ), 
            .Z(n30683));
    LUT4 mux_20_i86_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [85]), 
         .D(key_mem_new[85]), .Z(key_mem_0__127__N_5344[85])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i86_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25683 (.BLUT(n8_adj_9252), .ALUT(n9_adj_9251), .C0(\muxed_round_nr[1] ), 
          .Z(n30842));
    L6MUX21 i25525 (.D0(n30681), .D1(n33453), .SD(\muxed_round_nr[2] ), 
            .Z(n30684));
    LUT4 i3336_3_lut_4_lut (.A(prev_key1_reg[119]), .B(\round_key_gen.trw[23] ), 
         .C(n35835), .D(n33591), .Z(n8821)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam i3336_3_lut_4_lut.init = 16'hf606;
    L6MUX21 i25531 (.D0(n30686), .D1(n30687), .SD(\muxed_round_nr[2] ), 
            .Z(n30690));
    L6MUX21 i25532 (.D0(n30688), .D1(n33454), .SD(\muxed_round_nr[2] ), 
            .Z(n30691));
    LUT4 mux_20_i87_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [86]), 
         .D(key_mem_new[86]), .Z(key_mem_0__127__N_5344[86])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i87_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25688 (.BLUT(n1_adj_9249), .ALUT(n2_adj_9248), .C0(\muxed_round_nr[1] ), 
          .Z(n30847));
    LUT4 mux_51_i120_3_lut_4_lut (.A(prev_key1_reg[119]), .B(\round_key_gen.trw[23] ), 
         .C(n33860), .D(\key_reg[0] [23]), .Z(key_mem_new_127__N_7264[119])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam mux_51_i120_3_lut_4_lut.init = 16'h6f60;
    L6MUX21 i25538 (.D0(n30693), .D1(n30694), .SD(\muxed_round_nr[2] ), 
            .Z(n30697));
    LUT4 i3334_3_lut_4_lut (.A(prev_key1_reg[118]), .B(\round_key_gen.trw[22] ), 
         .C(n35835), .D(n33592), .Z(n8819)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam i3334_3_lut_4_lut.init = 16'hf606;
    L6MUX21 i25539 (.D0(n30695), .D1(n33455), .SD(\muxed_round_nr[2] ), 
            .Z(n30698));
    L6MUX21 i25545 (.D0(n30700), .D1(n30701), .SD(\muxed_round_nr[2] ), 
            .Z(n30704));
    PFUMX i25689 (.BLUT(n4_adj_9247), .ALUT(n5_adj_9246), .C0(\muxed_round_nr[1] ), 
          .Z(n30848));
    L6MUX21 i25546 (.D0(n30702), .D1(n33456), .SD(\muxed_round_nr[2] ), 
            .Z(n30705));
    L6MUX21 i25552 (.D0(n30707), .D1(n30708), .SD(\muxed_round_nr[2] ), 
            .Z(n30711));
    L6MUX21 i25553 (.D0(n30709), .D1(n33457), .SD(\muxed_round_nr[2] ), 
            .Z(n30712));
    LUT4 i11_4_lut_adj_658 (.A(n5), .B(keymem_sboxw[28]), .C(init_state), 
         .D(n10_adj_9264), .Z(muxed_sboxw[28])) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(181[17:28])
    defparam i11_4_lut_adj_658.init = 16'hc5c0;
    PFUMX i25690 (.BLUT(n8_adj_9245), .ALUT(n9_adj_9244), .C0(\muxed_round_nr[1] ), 
          .Z(n30849));
    L6MUX21 i25559 (.D0(n30714), .D1(n30715), .SD(\muxed_round_nr[2] ), 
            .Z(n30718));
    L6MUX21 i25560 (.D0(n30716), .D1(n33458), .SD(\muxed_round_nr[2] ), 
            .Z(n30719));
    LUT4 mux_51_i119_3_lut_4_lut (.A(prev_key1_reg[118]), .B(\round_key_gen.trw[22] ), 
         .C(n33860), .D(\key_reg[0] [22]), .Z(key_mem_new_127__N_7264[118])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam mux_51_i119_3_lut_4_lut.init = 16'h6f60;
    L6MUX21 i25566 (.D0(n30721), .D1(n30722), .SD(\muxed_round_nr[2] ), 
            .Z(n30725));
    L6MUX21 i25567 (.D0(n30723), .D1(n33459), .SD(\muxed_round_nr[2] ), 
            .Z(n30726));
    LUT4 mux_20_i88_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [87]), 
         .D(key_mem_new[87]), .Z(key_mem_0__127__N_5344[87])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i88_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i3332_3_lut_4_lut (.A(prev_key1_reg[117]), .B(\round_key_gen.trw[21] ), 
         .C(n35835), .D(n33593), .Z(n8817)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam i3332_3_lut_4_lut.init = 16'hf606;
    L6MUX21 i25573 (.D0(n30728), .D1(n30729), .SD(\muxed_round_nr[2] ), 
            .Z(n30732));
    LUT4 mux_85_i77_3_lut_rep_241_4_lut (.A(prev_key0_reg[76]), .B(n4_adj_8367), 
         .C(n33859), .D(\key_reg[5] [12]), .Z(n33545)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam mux_85_i77_3_lut_rep_241_4_lut.init = 16'h6f60;
    L6MUX21 i25574 (.D0(n30730), .D1(n33460), .SD(\muxed_round_nr[2] ), 
            .Z(n30733));
    PFUMX i25695 (.BLUT(n1_adj_9242), .ALUT(n2_adj_9241), .C0(\muxed_round_nr[1] ), 
          .Z(n30854));
    L6MUX21 i25580 (.D0(n30735), .D1(n30736), .SD(\muxed_round_nr[2] ), 
            .Z(n30739));
    L6MUX21 i25581 (.D0(n30737), .D1(n33461), .SD(\muxed_round_nr[2] ), 
            .Z(n30740));
    LUT4 round_3__I_0_Mux_102_i11_3_lut (.A(\key_mem[12] [102]), .B(\key_mem[13] [102]), 
         .C(n33952), .Z(n11_adj_124)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_102_i11_3_lut.init = 16'hcaca;
    PFUMX i25696 (.BLUT(n4_adj_9240), .ALUT(n5_adj_9239), .C0(\muxed_round_nr[1] ), 
          .Z(n30855));
    L6MUX21 i25587 (.D0(n30742), .D1(n30743), .SD(\muxed_round_nr[2] ), 
            .Z(n30746));
    L6MUX21 i25588 (.D0(n30744), .D1(n33462), .SD(\muxed_round_nr[2] ), 
            .Z(n30747));
    LUT4 mux_51_i118_3_lut_4_lut (.A(prev_key1_reg[117]), .B(\round_key_gen.trw[21] ), 
         .C(n33860), .D(\key_reg[0] [21]), .Z(key_mem_new_127__N_7264[117])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam mux_51_i118_3_lut_4_lut.init = 16'h6f60;
    LUT4 i3330_3_lut_4_lut (.A(prev_key1_reg[116]), .B(\round_key_gen.trw[20] ), 
         .C(n35835), .D(n33594), .Z(n8815)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam i3330_3_lut_4_lut.init = 16'hf606;
    L6MUX21 i25594 (.D0(n30749), .D1(n30750), .SD(\muxed_round_nr[2] ), 
            .Z(n30753));
    L6MUX21 i25595 (.D0(n30751), .D1(n33463), .SD(\muxed_round_nr[2] ), 
            .Z(n30754));
    LUT4 mux_51_i117_3_lut_4_lut (.A(prev_key1_reg[116]), .B(\round_key_gen.trw[20] ), 
         .C(n33860), .D(\key_reg[0] [20]), .Z(key_mem_new_127__N_7264[116])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam mux_51_i117_3_lut_4_lut.init = 16'h6f60;
    L6MUX21 i25601 (.D0(n30756), .D1(n30757), .SD(\muxed_round_nr[2] ), 
            .Z(n30760));
    L6MUX21 i25602 (.D0(n30758), .D1(n33336), .SD(\muxed_round_nr[2] ), 
            .Z(n30761));
    L6MUX21 i25608 (.D0(n30763), .D1(n30764), .SD(\muxed_round_nr[2] ), 
            .Z(n30767));
    PFUMX i25697 (.BLUT(n8_adj_9238), .ALUT(n9_adj_9237), .C0(\muxed_round_nr[1] ), 
          .Z(n30856));
    L6MUX21 i25609 (.D0(n30765), .D1(n33435), .SD(\muxed_round_nr[2] ), 
            .Z(n30768));
    L6MUX21 i25615 (.D0(n30770), .D1(n30771), .SD(\muxed_round_nr[2] ), 
            .Z(n30774));
    L6MUX21 i25616 (.D0(n30772), .D1(n33437), .SD(\muxed_round_nr[2] ), 
            .Z(n30775));
    LUT4 i3328_3_lut_4_lut (.A(prev_key1_reg[115]), .B(\round_key_gen.trw[19] ), 
         .C(n35835), .D(n33595), .Z(n8813)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam i3328_3_lut_4_lut.init = 16'hf606;
    LUT4 round_3__I_0_Mux_102_i9_3_lut (.A(\key_mem[10] [102]), .B(\key_mem[11] [102]), 
         .C(n33952), .Z(n9_adj_9266)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_102_i9_3_lut.init = 16'hcaca;
    L6MUX21 i25622 (.D0(n30777), .D1(n30778), .SD(\muxed_round_nr[2] ), 
            .Z(n30781));
    L6MUX21 i25623 (.D0(n30779), .D1(n33438), .SD(\muxed_round_nr[2] ), 
            .Z(n30782));
    LUT4 round_3__I_0_Mux_102_i8_3_lut (.A(\key_mem[8] [102]), .B(\key_mem[9] [102]), 
         .C(n33952), .Z(n8_adj_9267)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_102_i8_3_lut.init = 16'hcaca;
    LUT4 i11_4_lut_adj_659 (.A(n5), .B(keymem_sboxw[29]), .C(init_state), 
         .D(n10_adj_9268), .Z(muxed_sboxw[29])) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(181[17:28])
    defparam i11_4_lut_adj_659.init = 16'hc5c0;
    L6MUX21 i25629 (.D0(n30784), .D1(n30785), .SD(\muxed_round_nr[2] ), 
            .Z(n30788));
    L6MUX21 i25630 (.D0(n30786), .D1(n33439), .SD(\muxed_round_nr[2] ), 
            .Z(n30789));
    PFUMX i25702 (.BLUT(n1_adj_9235), .ALUT(n2_adj_9234), .C0(\muxed_round_nr[1] ), 
          .Z(n30861));
    LUT4 mux_51_i116_3_lut_4_lut (.A(prev_key1_reg[115]), .B(\round_key_gen.trw[19] ), 
         .C(n33860), .D(\key_reg[0] [19]), .Z(key_mem_new_127__N_7264[115])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam mux_51_i116_3_lut_4_lut.init = 16'h6f60;
    LUT4 i3326_3_lut_4_lut (.A(prev_key1_reg[114]), .B(\round_key_gen.trw[18] ), 
         .C(n35835), .D(n33596), .Z(n8811)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam i3326_3_lut_4_lut.init = 16'hf606;
    L6MUX21 i25636 (.D0(n30791), .D1(n30792), .SD(\muxed_round_nr[2] ), 
            .Z(n30795));
    L6MUX21 i25637 (.D0(n30793), .D1(n33440), .SD(\muxed_round_nr[2] ), 
            .Z(n30796));
    LUT4 mux_51_i115_3_lut_4_lut (.A(prev_key1_reg[114]), .B(\round_key_gen.trw[18] ), 
         .C(n33860), .D(\key_reg[0] [18]), .Z(key_mem_new_127__N_7264[114])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam mux_51_i115_3_lut_4_lut.init = 16'h6f60;
    PFUMX i25703 (.BLUT(n4_adj_9233), .ALUT(n5_adj_9232), .C0(\muxed_round_nr[1] ), 
          .Z(n30862));
    L6MUX21 i25643 (.D0(n30798), .D1(n30799), .SD(\muxed_round_nr[2] ), 
            .Z(n30802));
    L6MUX21 i25644 (.D0(n30800), .D1(n33442), .SD(\muxed_round_nr[2] ), 
            .Z(n30803));
    PFUMX i25704 (.BLUT(n8_adj_9231), .ALUT(n9_adj_9230), .C0(\muxed_round_nr[1] ), 
          .Z(n30863));
    LUT4 i3324_3_lut_4_lut (.A(prev_key1_reg[113]), .B(\round_key_gen.trw[17] ), 
         .C(n35835), .D(n33597), .Z(n8809)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam i3324_3_lut_4_lut.init = 16'hf606;
    L6MUX21 i25650 (.D0(n30805), .D1(n30806), .SD(\muxed_round_nr[2] ), 
            .Z(n30809));
    LUT4 mux_20_i89_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [88]), 
         .D(key_mem_new[88]), .Z(key_mem_0__127__N_5344[88])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i89_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i90_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [89]), 
         .D(key_mem_new[89]), .Z(key_mem_0__127__N_5344[89])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i90_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i91_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [90]), 
         .D(key_mem_new[90]), .Z(key_mem_0__127__N_5344[90])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i91_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i92_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [91]), 
         .D(key_mem_new[91]), .Z(key_mem_0__127__N_5344[91])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i92_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i93_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [92]), 
         .D(key_mem_new[92]), .Z(key_mem_0__127__N_5344[92])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i93_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i94_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [93]), 
         .D(key_mem_new[93]), .Z(key_mem_0__127__N_5344[93])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i94_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i95_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [94]), 
         .D(key_mem_new[94]), .Z(key_mem_0__127__N_5344[94])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i95_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i96_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [95]), 
         .D(key_mem_new[95]), .Z(key_mem_0__127__N_5344[95])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i96_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i97_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [96]), 
         .D(key_mem_new[96]), .Z(key_mem_0__127__N_5344[96])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i97_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i98_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [97]), 
         .D(key_mem_new[97]), .Z(key_mem_0__127__N_5344[97])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i98_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i99_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [98]), 
         .D(key_mem_new[98]), .Z(key_mem_0__127__N_5344[98])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i99_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i100_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [99]), 
         .D(key_mem_new[99]), .Z(key_mem_0__127__N_5344[99])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i100_3_lut_4_lut.init = 16'hf2d0;
    LUT4 round_3__I_0_Mux_102_i5_3_lut (.A(\key_mem[6] [102]), .B(\key_mem[7] [102]), 
         .C(n33952), .Z(n5_adj_9269)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_102_i5_3_lut.init = 16'hcaca;
    L6MUX21 i25651 (.D0(n30807), .D1(n33443), .SD(\muxed_round_nr[2] ), 
            .Z(n30810));
    L6MUX21 i25657 (.D0(n30812), .D1(n30813), .SD(\muxed_round_nr[2] ), 
            .Z(n30816));
    LUT4 i11_4_lut_adj_660 (.A(n5), .B(keymem_sboxw[30]), .C(init_state), 
         .D(n10_adj_9270), .Z(muxed_sboxw[30])) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(181[17:28])
    defparam i11_4_lut_adj_660.init = 16'hc5c0;
    L6MUX21 i25658 (.D0(n30814), .D1(n33444), .SD(\muxed_round_nr[2] ), 
            .Z(n30817));
    LUT4 round_3__I_0_Mux_102_i4_3_lut (.A(\key_mem[4] [102]), .B(\key_mem[5] [102]), 
         .C(n33952), .Z(n4_adj_9271)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_102_i4_3_lut.init = 16'hcaca;
    LUT4 mux_51_i114_3_lut_4_lut (.A(prev_key1_reg[113]), .B(\round_key_gen.trw[17] ), 
         .C(n33860), .D(\key_reg[0] [17]), .Z(key_mem_new_127__N_7264[113])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam mux_51_i114_3_lut_4_lut.init = 16'h6f60;
    LUT4 i11_4_lut_adj_661 (.A(n5), .B(keymem_sboxw[31]), .C(init_state), 
         .D(n10_adj_9272), .Z(muxed_sboxw[31])) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(181[17:28])
    defparam i11_4_lut_adj_661.init = 16'hc5c0;
    L6MUX21 i25664 (.D0(n30819), .D1(n30820), .SD(\muxed_round_nr[2] ), 
            .Z(n30823));
    L6MUX21 i25665 (.D0(n30821), .D1(n33445), .SD(\muxed_round_nr[2] ), 
            .Z(n30824));
    L6MUX21 i25671 (.D0(n30826), .D1(n30827), .SD(\muxed_round_nr[2] ), 
            .Z(n30830));
    L6MUX21 i25672 (.D0(n30828), .D1(n33447), .SD(\muxed_round_nr[2] ), 
            .Z(n30831));
    PFUMX i25709 (.BLUT(n1_adj_9228), .ALUT(n2_adj_9227), .C0(\muxed_round_nr[1] ), 
          .Z(n30868));
    L6MUX21 i25678 (.D0(n30833), .D1(n30834), .SD(\muxed_round_nr[2] ), 
            .Z(n30837));
    LUT4 i3322_3_lut_4_lut (.A(prev_key1_reg[112]), .B(\round_key_gen.trw[16] ), 
         .C(n35835), .D(n33598), .Z(n8807)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam i3322_3_lut_4_lut.init = 16'hf606;
    L6MUX21 i25679 (.D0(n30835), .D1(n33337), .SD(\muxed_round_nr[2] ), 
            .Z(n30838));
    LUT4 mux_20_i101_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [100]), 
         .D(key_mem_new[100]), .Z(key_mem_0__127__N_5344[100])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i101_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25710 (.BLUT(n4_adj_9226), .ALUT(n5_adj_9225), .C0(\muxed_round_nr[1] ), 
          .Z(n30869));
    L6MUX21 i25685 (.D0(n30840), .D1(n30841), .SD(\muxed_round_nr[2] ), 
            .Z(n30844));
    LUT4 round_3__I_0_Mux_102_i2_3_lut (.A(\key_mem[2] [102]), .B(\key_mem[3] [102]), 
         .C(n33952), .Z(n2_adj_9273)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_102_i2_3_lut.init = 16'hcaca;
    L6MUX21 i25686 (.D0(n30842), .D1(n33338), .SD(\muxed_round_nr[2] ), 
            .Z(n30845));
    L6MUX21 i25692 (.D0(n30847), .D1(n30848), .SD(\muxed_round_nr[2] ), 
            .Z(n30851));
    L6MUX21 i25693 (.D0(n30849), .D1(n33339), .SD(\muxed_round_nr[2] ), 
            .Z(n30852));
    L6MUX21 i25699 (.D0(n30854), .D1(n30855), .SD(\muxed_round_nr[2] ), 
            .Z(n30858));
    PFUMX i25711 (.BLUT(n8_adj_9224), .ALUT(n9_adj_9223), .C0(\muxed_round_nr[1] ), 
          .Z(n30870));
    L6MUX21 i25700 (.D0(n30856), .D1(n33340), .SD(\muxed_round_nr[2] ), 
            .Z(n30859));
    L6MUX21 i25706 (.D0(n30861), .D1(n30862), .SD(\muxed_round_nr[2] ), 
            .Z(n30865));
    LUT4 mux_51_i113_3_lut_4_lut (.A(prev_key1_reg[112]), .B(\round_key_gen.trw[16] ), 
         .C(n33860), .D(\key_reg[0] [16]), .Z(key_mem_new_127__N_7264[112])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam mux_51_i113_3_lut_4_lut.init = 16'h6f60;
    LUT4 i3320_3_lut_4_lut (.A(prev_key1_reg[111]), .B(\round_key_gen.trw[15] ), 
         .C(n35835), .D(n33599), .Z(n8805)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam i3320_3_lut_4_lut.init = 16'hf606;
    L6MUX21 i25707 (.D0(n30863), .D1(n33341), .SD(\muxed_round_nr[2] ), 
            .Z(n30866));
    L6MUX21 i25713 (.D0(n30868), .D1(n30869), .SD(\muxed_round_nr[2] ), 
            .Z(n30872));
    LUT4 mux_20_i102_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [101]), 
         .D(key_mem_new[101]), .Z(key_mem_0__127__N_5344[101])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i102_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i103_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [102]), 
         .D(key_mem_new[102]), .Z(key_mem_0__127__N_5344[102])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i103_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i104_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [103]), 
         .D(key_mem_new[103]), .Z(key_mem_0__127__N_5344[103])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i104_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i105_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [104]), 
         .D(key_mem_new[104]), .Z(key_mem_0__127__N_5344[104])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i105_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i106_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [105]), 
         .D(key_mem_new[105]), .Z(key_mem_0__127__N_5344[105])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i106_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i107_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [106]), 
         .D(key_mem_new[106]), .Z(key_mem_0__127__N_5344[106])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i107_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i108_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [107]), 
         .D(key_mem_new[107]), .Z(key_mem_0__127__N_5344[107])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i108_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i109_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [108]), 
         .D(key_mem_new[108]), .Z(key_mem_0__127__N_5344[108])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i109_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i110_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [109]), 
         .D(key_mem_new[109]), .Z(key_mem_0__127__N_5344[109])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i110_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i111_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [110]), 
         .D(key_mem_new[110]), .Z(key_mem_0__127__N_5344[110])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i111_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i112_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [111]), 
         .D(key_mem_new[111]), .Z(key_mem_0__127__N_5344[111])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i112_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i113_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [112]), 
         .D(key_mem_new[112]), .Z(key_mem_0__127__N_5344[112])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i113_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i114_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [113]), 
         .D(key_mem_new[113]), .Z(key_mem_0__127__N_5344[113])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i114_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i115_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [114]), 
         .D(key_mem_new[114]), .Z(key_mem_0__127__N_5344[114])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i115_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i116_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [115]), 
         .D(key_mem_new[115]), .Z(key_mem_0__127__N_5344[115])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i116_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i117_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [116]), 
         .D(key_mem_new[116]), .Z(key_mem_0__127__N_5344[116])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i117_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i118_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [117]), 
         .D(key_mem_new[117]), .Z(key_mem_0__127__N_5344[117])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i118_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i119_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [118]), 
         .D(key_mem_new[118]), .Z(key_mem_0__127__N_5344[118])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i119_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i120_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [119]), 
         .D(key_mem_new[119]), .Z(key_mem_0__127__N_5344[119])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i120_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i121_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [120]), 
         .D(key_mem_new[120]), .Z(key_mem_0__127__N_5344[120])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i121_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i122_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [121]), 
         .D(key_mem_new[121]), .Z(key_mem_0__127__N_5344[121])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i122_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i123_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [122]), 
         .D(key_mem_new[122]), .Z(key_mem_0__127__N_5344[122])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i123_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i124_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [123]), 
         .D(key_mem_new[123]), .Z(key_mem_0__127__N_5344[123])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i124_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i125_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [124]), 
         .D(key_mem_new[124]), .Z(key_mem_0__127__N_5344[124])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i125_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i126_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [125]), 
         .D(key_mem_new[125]), .Z(key_mem_0__127__N_5344[125])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i126_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i127_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [126]), 
         .D(key_mem_new[126]), .Z(key_mem_0__127__N_5344[126])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i127_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i128_3_lut_4_lut (.A(n33938), .B(n33944), .C(\key_mem[3] [127]), 
         .D(key_mem_new[127]), .Z(key_mem_0__127__N_5344[127])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_20_i128_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_19_i1_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [0]), 
         .D(key_mem_new[0]), .Z(key_mem_0__127__N_5472[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i2_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [1]), 
         .D(key_mem_new[1]), .Z(key_mem_0__127__N_5472[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i3_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [2]), 
         .D(key_mem_new[2]), .Z(key_mem_0__127__N_5472[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i4_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [3]), 
         .D(key_mem_new[3]), .Z(key_mem_0__127__N_5472[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i5_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [4]), 
         .D(key_mem_new[4]), .Z(key_mem_0__127__N_5472[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i6_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [5]), 
         .D(key_mem_new[5]), .Z(key_mem_0__127__N_5472[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i7_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [6]), 
         .D(key_mem_new[6]), .Z(key_mem_0__127__N_5472[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i8_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [7]), 
         .D(key_mem_new[7]), .Z(key_mem_0__127__N_5472[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i9_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [8]), 
         .D(key_mem_new[8]), .Z(key_mem_0__127__N_5472[8])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i9_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i10_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [9]), 
         .D(key_mem_new[9]), .Z(key_mem_0__127__N_5472[9])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i10_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i11_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [10]), 
         .D(key_mem_new[10]), .Z(key_mem_0__127__N_5472[10])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i11_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i12_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [11]), 
         .D(key_mem_new[11]), .Z(key_mem_0__127__N_5472[11])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i12_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i13_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [12]), 
         .D(key_mem_new[12]), .Z(key_mem_0__127__N_5472[12])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i13_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i14_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [13]), 
         .D(key_mem_new[13]), .Z(key_mem_0__127__N_5472[13])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i14_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i15_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [14]), 
         .D(key_mem_new[14]), .Z(key_mem_0__127__N_5472[14])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i15_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i16_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [15]), 
         .D(key_mem_new[15]), .Z(key_mem_0__127__N_5472[15])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i16_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i17_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [16]), 
         .D(key_mem_new[16]), .Z(key_mem_0__127__N_5472[16])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i17_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i18_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [17]), 
         .D(key_mem_new[17]), .Z(key_mem_0__127__N_5472[17])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i18_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i19_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [18]), 
         .D(key_mem_new[18]), .Z(key_mem_0__127__N_5472[18])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i19_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i20_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [19]), 
         .D(key_mem_new[19]), .Z(key_mem_0__127__N_5472[19])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i20_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i21_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [20]), 
         .D(key_mem_new[20]), .Z(key_mem_0__127__N_5472[20])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i21_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i22_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [21]), 
         .D(key_mem_new[21]), .Z(key_mem_0__127__N_5472[21])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i22_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i23_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [22]), 
         .D(key_mem_new[22]), .Z(key_mem_0__127__N_5472[22])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i23_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i24_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [23]), 
         .D(key_mem_new[23]), .Z(key_mem_0__127__N_5472[23])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i24_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i25_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [24]), 
         .D(key_mem_new[24]), .Z(key_mem_0__127__N_5472[24])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i25_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i26_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [25]), 
         .D(key_mem_new[25]), .Z(key_mem_0__127__N_5472[25])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i26_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i27_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [26]), 
         .D(key_mem_new[26]), .Z(key_mem_0__127__N_5472[26])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i27_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i28_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [27]), 
         .D(key_mem_new[27]), .Z(key_mem_0__127__N_5472[27])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i28_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i29_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [28]), 
         .D(key_mem_new[28]), .Z(key_mem_0__127__N_5472[28])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i29_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i30_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [29]), 
         .D(key_mem_new[29]), .Z(key_mem_0__127__N_5472[29])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i30_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i31_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [30]), 
         .D(key_mem_new[30]), .Z(key_mem_0__127__N_5472[30])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i31_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i32_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [31]), 
         .D(key_mem_new[31]), .Z(key_mem_0__127__N_5472[31])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i32_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i33_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [32]), 
         .D(key_mem_new[32]), .Z(key_mem_0__127__N_5472[32])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i33_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i34_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [33]), 
         .D(key_mem_new[33]), .Z(key_mem_0__127__N_5472[33])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i34_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i35_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [34]), 
         .D(key_mem_new[34]), .Z(key_mem_0__127__N_5472[34])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i35_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i36_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [35]), 
         .D(key_mem_new[35]), .Z(key_mem_0__127__N_5472[35])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i36_3_lut_4_lut.init = 16'hf1e0;
    L6MUX21 i25714 (.D0(n30870), .D1(n33342), .SD(\muxed_round_nr[2] ), 
            .Z(n30873));
    LUT4 round_3__I_0_Mux_102_i1_3_lut (.A(\key_mem[0] [102]), .B(\key_mem[1] [102]), 
         .C(n33952), .Z(n1_adj_9274)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_102_i1_3_lut.init = 16'hcaca;
    LUT4 mux_19_i37_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [36]), 
         .D(key_mem_new[36]), .Z(key_mem_0__127__N_5472[36])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i37_3_lut_4_lut.init = 16'hf1e0;
    L6MUX21 i25720 (.D0(n30875), .D1(n30876), .SD(\muxed_round_nr[2] ), 
            .Z(n30879));
    PFUMX i25716 (.BLUT(n1_adj_9221), .ALUT(n2_adj_9220), .C0(\muxed_round_nr[1] ), 
          .Z(n30875));
    L6MUX21 i25721 (.D0(n30877), .D1(n33350), .SD(\muxed_round_nr[2] ), 
            .Z(n30880));
    LUT4 mux_51_i112_3_lut_4_lut (.A(prev_key1_reg[111]), .B(\round_key_gen.trw[15] ), 
         .C(n33860), .D(\key_reg[0] [15]), .Z(key_mem_new_127__N_7264[111])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam mux_51_i112_3_lut_4_lut.init = 16'h6f60;
    LUT4 i3318_3_lut_4_lut (.A(prev_key1_reg[110]), .B(\round_key_gen.trw[14] ), 
         .C(n35835), .D(n33600), .Z(n8803)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam i3318_3_lut_4_lut.init = 16'hf606;
    L6MUX21 i25727 (.D0(n30882), .D1(n30883), .SD(\muxed_round_nr[2] ), 
            .Z(n30886));
    L6MUX21 i25728 (.D0(n30884), .D1(n33355), .SD(\muxed_round_nr[2] ), 
            .Z(n30887));
    PFUMX i25717 (.BLUT(n4_adj_9216), .ALUT(n5_adj_9215), .C0(\muxed_round_nr[1] ), 
          .Z(n30876));
    LUT4 i6_2_lut_3_lut_adj_662 (.A(prev_key1_reg[43]), .B(n33736), .C(keymem_sboxw[11]), 
         .Z(n16017)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;
    defparam i6_2_lut_3_lut_adj_662.init = 16'h9696;
    LUT4 mux_51_i111_3_lut_4_lut (.A(prev_key1_reg[110]), .B(\round_key_gen.trw[14] ), 
         .C(n33860), .D(\key_reg[0] [14]), .Z(key_mem_new_127__N_7264[110])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam mux_51_i111_3_lut_4_lut.init = 16'h6f60;
    L6MUX21 i25734 (.D0(n30889), .D1(n30890), .SD(\muxed_round_nr[2] ), 
            .Z(n30893));
    L6MUX21 i25735 (.D0(n30891), .D1(n33361), .SD(\muxed_round_nr[2] ), 
            .Z(n30894));
    L6MUX21 i25741 (.D0(n30896), .D1(n30897), .SD(\muxed_round_nr[2] ), 
            .Z(n30900));
    L6MUX21 i25742 (.D0(n30898), .D1(n33367), .SD(\muxed_round_nr[2] ), 
            .Z(n30901));
    LUT4 i3316_3_lut_4_lut (.A(prev_key1_reg[109]), .B(\round_key_gen.trw[13] ), 
         .C(n35835), .D(n33601), .Z(n8801)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam i3316_3_lut_4_lut.init = 16'hf606;
    L6MUX21 i25748 (.D0(n30903), .D1(n30904), .SD(\muxed_round_nr[2] ), 
            .Z(n30907));
    L6MUX21 i25749 (.D0(n30905), .D1(n33374), .SD(\muxed_round_nr[2] ), 
            .Z(n30908));
    LUT4 mux_51_i110_3_lut_4_lut (.A(prev_key1_reg[109]), .B(\round_key_gen.trw[13] ), 
         .C(n33860), .D(\key_reg[0] [13]), .Z(key_mem_new_127__N_7264[109])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam mux_51_i110_3_lut_4_lut.init = 16'h6f60;
    L6MUX21 i25755 (.D0(n30910), .D1(n30911), .SD(\muxed_round_nr[2] ), 
            .Z(n30914));
    L6MUX21 i25756 (.D0(n30912), .D1(n33377), .SD(\muxed_round_nr[2] ), 
            .Z(n30915));
    LUT4 mux_19_i38_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [37]), 
         .D(key_mem_new[37]), .Z(key_mem_0__127__N_5472[37])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i38_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i39_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [38]), 
         .D(key_mem_new[38]), .Z(key_mem_0__127__N_5472[38])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i39_3_lut_4_lut.init = 16'hf1e0;
    L6MUX21 i25762 (.D0(n30917), .D1(n30918), .SD(\muxed_round_nr[2] ), 
            .Z(n30921));
    L6MUX21 i25763 (.D0(n30919), .D1(n33379), .SD(\muxed_round_nr[2] ), 
            .Z(n30922));
    L6MUX21 i25865 (.D0(n31020), .D1(n31021), .SD(\muxed_round_nr[2] ), 
            .Z(n31024));
    LUT4 i3314_3_lut_4_lut (.A(prev_key1_reg[108]), .B(\round_key_gen.trw[12] ), 
         .C(n35835), .D(n33602), .Z(n8799)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam i3314_3_lut_4_lut.init = 16'hf606;
    L6MUX21 i25866 (.D0(n31022), .D1(n33380), .SD(\muxed_round_nr[2] ), 
            .Z(n31025));
    L6MUX21 i25872 (.D0(n31027), .D1(n31028), .SD(\muxed_round_nr[2] ), 
            .Z(n31031));
    LUT4 mux_19_i40_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [39]), 
         .D(key_mem_new[39]), .Z(key_mem_0__127__N_5472[39])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i40_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i41_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [40]), 
         .D(key_mem_new[40]), .Z(key_mem_0__127__N_5472[40])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i41_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i42_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [41]), 
         .D(key_mem_new[41]), .Z(key_mem_0__127__N_5472[41])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i42_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i43_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [42]), 
         .D(key_mem_new[42]), .Z(key_mem_0__127__N_5472[42])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i43_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i44_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [43]), 
         .D(key_mem_new[43]), .Z(key_mem_0__127__N_5472[43])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i44_3_lut_4_lut.init = 16'hf1e0;
    L6MUX21 i25873 (.D0(n31029), .D1(n33382), .SD(\muxed_round_nr[2] ), 
            .Z(n31032));
    LUT4 mux_19_i45_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [44]), 
         .D(key_mem_new[44]), .Z(key_mem_0__127__N_5472[44])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i45_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i46_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [45]), 
         .D(key_mem_new[45]), .Z(key_mem_0__127__N_5472[45])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i46_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_51_i109_3_lut_4_lut (.A(prev_key1_reg[108]), .B(\round_key_gen.trw[12] ), 
         .C(n33860), .D(\key_reg[0] [12]), .Z(key_mem_new_127__N_7264[108])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam mux_51_i109_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_19_i47_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [46]), 
         .D(key_mem_new[46]), .Z(key_mem_0__127__N_5472[46])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i47_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3312_3_lut_4_lut (.A(prev_key1_reg[107]), .B(\round_key_gen.trw[11] ), 
         .C(n35835), .D(n33603), .Z(n8797)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam i3312_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_19_i48_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [47]), 
         .D(key_mem_new[47]), .Z(key_mem_0__127__N_5472[47])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i48_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i49_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [48]), 
         .D(key_mem_new[48]), .Z(key_mem_0__127__N_5472[48])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i49_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i50_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [49]), 
         .D(key_mem_new[49]), .Z(key_mem_0__127__N_5472[49])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i50_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i51_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [50]), 
         .D(key_mem_new[50]), .Z(key_mem_0__127__N_5472[50])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i51_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i52_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [51]), 
         .D(key_mem_new[51]), .Z(key_mem_0__127__N_5472[51])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i52_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i53_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [52]), 
         .D(key_mem_new[52]), .Z(key_mem_0__127__N_5472[52])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i53_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i54_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [53]), 
         .D(key_mem_new[53]), .Z(key_mem_0__127__N_5472[53])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i54_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i55_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [54]), 
         .D(key_mem_new[54]), .Z(key_mem_0__127__N_5472[54])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i55_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i56_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [55]), 
         .D(key_mem_new[55]), .Z(key_mem_0__127__N_5472[55])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i56_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i57_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [56]), 
         .D(key_mem_new[56]), .Z(key_mem_0__127__N_5472[56])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i57_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i58_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [57]), 
         .D(key_mem_new[57]), .Z(key_mem_0__127__N_5472[57])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i58_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i59_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [58]), 
         .D(key_mem_new[58]), .Z(key_mem_0__127__N_5472[58])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i59_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i60_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [59]), 
         .D(key_mem_new[59]), .Z(key_mem_0__127__N_5472[59])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i60_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i61_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [60]), 
         .D(key_mem_new[60]), .Z(key_mem_0__127__N_5472[60])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i61_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i62_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [61]), 
         .D(key_mem_new[61]), .Z(key_mem_0__127__N_5472[61])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i62_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i63_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [62]), 
         .D(key_mem_new[62]), .Z(key_mem_0__127__N_5472[62])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i63_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i64_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [63]), 
         .D(key_mem_new[63]), .Z(key_mem_0__127__N_5472[63])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i64_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i65_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [64]), 
         .D(key_mem_new[64]), .Z(key_mem_0__127__N_5472[64])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i65_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i66_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [65]), 
         .D(key_mem_new[65]), .Z(key_mem_0__127__N_5472[65])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i66_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i67_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [66]), 
         .D(key_mem_new[66]), .Z(key_mem_0__127__N_5472[66])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i67_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i68_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [67]), 
         .D(key_mem_new[67]), .Z(key_mem_0__127__N_5472[67])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i68_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i69_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [68]), 
         .D(key_mem_new[68]), .Z(key_mem_0__127__N_5472[68])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i69_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i70_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [69]), 
         .D(key_mem_new[69]), .Z(key_mem_0__127__N_5472[69])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i70_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i71_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [70]), 
         .D(key_mem_new[70]), .Z(key_mem_0__127__N_5472[70])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i71_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i72_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [71]), 
         .D(key_mem_new[71]), .Z(key_mem_0__127__N_5472[71])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i72_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i73_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [72]), 
         .D(key_mem_new[72]), .Z(key_mem_0__127__N_5472[72])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i73_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i74_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [73]), 
         .D(key_mem_new[73]), .Z(key_mem_0__127__N_5472[73])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i74_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i75_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [74]), 
         .D(key_mem_new[74]), .Z(key_mem_0__127__N_5472[74])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i75_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i76_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [75]), 
         .D(key_mem_new[75]), .Z(key_mem_0__127__N_5472[75])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i76_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i77_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [76]), 
         .D(key_mem_new[76]), .Z(key_mem_0__127__N_5472[76])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i77_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i78_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [77]), 
         .D(key_mem_new[77]), .Z(key_mem_0__127__N_5472[77])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i78_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i79_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [78]), 
         .D(key_mem_new[78]), .Z(key_mem_0__127__N_5472[78])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i79_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i80_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [79]), 
         .D(key_mem_new[79]), .Z(key_mem_0__127__N_5472[79])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i80_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i81_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [80]), 
         .D(key_mem_new[80]), .Z(key_mem_0__127__N_5472[80])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i81_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i82_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [81]), 
         .D(key_mem_new[81]), .Z(key_mem_0__127__N_5472[81])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i82_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i83_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [82]), 
         .D(key_mem_new[82]), .Z(key_mem_0__127__N_5472[82])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i83_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i84_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [83]), 
         .D(key_mem_new[83]), .Z(key_mem_0__127__N_5472[83])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i84_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i85_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [84]), 
         .D(key_mem_new[84]), .Z(key_mem_0__127__N_5472[84])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i85_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i86_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [85]), 
         .D(key_mem_new[85]), .Z(key_mem_0__127__N_5472[85])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i86_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i87_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [86]), 
         .D(key_mem_new[86]), .Z(key_mem_0__127__N_5472[86])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i87_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i88_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [87]), 
         .D(key_mem_new[87]), .Z(key_mem_0__127__N_5472[87])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i88_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i89_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [88]), 
         .D(key_mem_new[88]), .Z(key_mem_0__127__N_5472[88])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i89_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i90_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [89]), 
         .D(key_mem_new[89]), .Z(key_mem_0__127__N_5472[89])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i90_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i91_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [90]), 
         .D(key_mem_new[90]), .Z(key_mem_0__127__N_5472[90])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i91_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i92_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [91]), 
         .D(key_mem_new[91]), .Z(key_mem_0__127__N_5472[91])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i92_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i93_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [92]), 
         .D(key_mem_new[92]), .Z(key_mem_0__127__N_5472[92])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i93_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i94_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [93]), 
         .D(key_mem_new[93]), .Z(key_mem_0__127__N_5472[93])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i94_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i95_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [94]), 
         .D(key_mem_new[94]), .Z(key_mem_0__127__N_5472[94])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i95_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i96_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [95]), 
         .D(key_mem_new[95]), .Z(key_mem_0__127__N_5472[95])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i96_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i97_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [96]), 
         .D(key_mem_new[96]), .Z(key_mem_0__127__N_5472[96])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i97_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i98_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [97]), 
         .D(key_mem_new[97]), .Z(key_mem_0__127__N_5472[97])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i98_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i99_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [98]), 
         .D(key_mem_new[98]), .Z(key_mem_0__127__N_5472[98])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i99_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i100_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [99]), 
         .D(key_mem_new[99]), .Z(key_mem_0__127__N_5472[99])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i100_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i101_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [100]), 
         .D(key_mem_new[100]), .Z(key_mem_0__127__N_5472[100])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i101_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i102_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [101]), 
         .D(key_mem_new[101]), .Z(key_mem_0__127__N_5472[101])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i102_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i103_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [102]), 
         .D(key_mem_new[102]), .Z(key_mem_0__127__N_5472[102])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i103_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i104_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [103]), 
         .D(key_mem_new[103]), .Z(key_mem_0__127__N_5472[103])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i104_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i105_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [104]), 
         .D(key_mem_new[104]), .Z(key_mem_0__127__N_5472[104])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i105_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i106_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [105]), 
         .D(key_mem_new[105]), .Z(key_mem_0__127__N_5472[105])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i106_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i107_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [106]), 
         .D(key_mem_new[106]), .Z(key_mem_0__127__N_5472[106])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i107_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i108_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [107]), 
         .D(key_mem_new[107]), .Z(key_mem_0__127__N_5472[107])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i108_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i109_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [108]), 
         .D(key_mem_new[108]), .Z(key_mem_0__127__N_5472[108])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i109_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i110_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [109]), 
         .D(key_mem_new[109]), .Z(key_mem_0__127__N_5472[109])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i110_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i111_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [110]), 
         .D(key_mem_new[110]), .Z(key_mem_0__127__N_5472[110])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i111_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i112_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [111]), 
         .D(key_mem_new[111]), .Z(key_mem_0__127__N_5472[111])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i112_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i113_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [112]), 
         .D(key_mem_new[112]), .Z(key_mem_0__127__N_5472[112])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i113_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i114_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [113]), 
         .D(key_mem_new[113]), .Z(key_mem_0__127__N_5472[113])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i114_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i115_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [114]), 
         .D(key_mem_new[114]), .Z(key_mem_0__127__N_5472[114])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i115_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i116_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [115]), 
         .D(key_mem_new[115]), .Z(key_mem_0__127__N_5472[115])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i116_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i117_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [116]), 
         .D(key_mem_new[116]), .Z(key_mem_0__127__N_5472[116])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i117_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i118_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [117]), 
         .D(key_mem_new[117]), .Z(key_mem_0__127__N_5472[117])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i118_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i119_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [118]), 
         .D(key_mem_new[118]), .Z(key_mem_0__127__N_5472[118])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i119_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i120_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [119]), 
         .D(key_mem_new[119]), .Z(key_mem_0__127__N_5472[119])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i120_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i121_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [120]), 
         .D(key_mem_new[120]), .Z(key_mem_0__127__N_5472[120])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i121_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i122_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [121]), 
         .D(key_mem_new[121]), .Z(key_mem_0__127__N_5472[121])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i122_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i123_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [122]), 
         .D(key_mem_new[122]), .Z(key_mem_0__127__N_5472[122])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i123_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i124_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [123]), 
         .D(key_mem_new[123]), .Z(key_mem_0__127__N_5472[123])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i124_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i125_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [124]), 
         .D(key_mem_new[124]), .Z(key_mem_0__127__N_5472[124])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i125_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i126_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [125]), 
         .D(key_mem_new[125]), .Z(key_mem_0__127__N_5472[125])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i126_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i127_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [126]), 
         .D(key_mem_new[126]), .Z(key_mem_0__127__N_5472[126])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i127_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19_i128_3_lut_4_lut (.A(n33943), .B(n33916), .C(\key_mem[4] [127]), 
         .D(key_mem_new[127]), .Z(key_mem_0__127__N_5472[127])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_19_i128_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i1_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [0]), 
         .D(key_mem_new[0]), .Z(key_mem_0__127__N_5600[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i2_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [1]), 
         .D(key_mem_new[1]), .Z(key_mem_0__127__N_5600[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i3_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [2]), 
         .D(key_mem_new[2]), .Z(key_mem_0__127__N_5600[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i4_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [3]), 
         .D(key_mem_new[3]), .Z(key_mem_0__127__N_5600[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i5_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [4]), 
         .D(key_mem_new[4]), .Z(key_mem_0__127__N_5600[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i6_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [5]), 
         .D(key_mem_new[5]), .Z(key_mem_0__127__N_5600[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i7_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [6]), 
         .D(key_mem_new[6]), .Z(key_mem_0__127__N_5600[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i8_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [7]), 
         .D(key_mem_new[7]), .Z(key_mem_0__127__N_5600[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i9_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [8]), 
         .D(key_mem_new[8]), .Z(key_mem_0__127__N_5600[8])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i9_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i10_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [9]), 
         .D(key_mem_new[9]), .Z(key_mem_0__127__N_5600[9])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i10_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i11_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [10]), 
         .D(key_mem_new[10]), .Z(key_mem_0__127__N_5600[10])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i11_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i12_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [11]), 
         .D(key_mem_new[11]), .Z(key_mem_0__127__N_5600[11])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i12_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i13_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [12]), 
         .D(key_mem_new[12]), .Z(key_mem_0__127__N_5600[12])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i13_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i14_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [13]), 
         .D(key_mem_new[13]), .Z(key_mem_0__127__N_5600[13])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i14_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i15_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [14]), 
         .D(key_mem_new[14]), .Z(key_mem_0__127__N_5600[14])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i15_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i16_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [15]), 
         .D(key_mem_new[15]), .Z(key_mem_0__127__N_5600[15])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i16_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i17_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [16]), 
         .D(key_mem_new[16]), .Z(key_mem_0__127__N_5600[16])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i17_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i18_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [17]), 
         .D(key_mem_new[17]), .Z(key_mem_0__127__N_5600[17])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i18_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i19_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [18]), 
         .D(key_mem_new[18]), .Z(key_mem_0__127__N_5600[18])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i19_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i20_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [19]), 
         .D(key_mem_new[19]), .Z(key_mem_0__127__N_5600[19])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i20_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i21_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [20]), 
         .D(key_mem_new[20]), .Z(key_mem_0__127__N_5600[20])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i21_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i22_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [21]), 
         .D(key_mem_new[21]), .Z(key_mem_0__127__N_5600[21])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i22_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i23_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [22]), 
         .D(key_mem_new[22]), .Z(key_mem_0__127__N_5600[22])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i23_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i24_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [23]), 
         .D(key_mem_new[23]), .Z(key_mem_0__127__N_5600[23])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i24_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i25_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [24]), 
         .D(key_mem_new[24]), .Z(key_mem_0__127__N_5600[24])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i25_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i26_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [25]), 
         .D(key_mem_new[25]), .Z(key_mem_0__127__N_5600[25])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i26_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i27_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [26]), 
         .D(key_mem_new[26]), .Z(key_mem_0__127__N_5600[26])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i27_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i28_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [27]), 
         .D(key_mem_new[27]), .Z(key_mem_0__127__N_5600[27])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i28_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i29_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [28]), 
         .D(key_mem_new[28]), .Z(key_mem_0__127__N_5600[28])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i29_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i30_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [29]), 
         .D(key_mem_new[29]), .Z(key_mem_0__127__N_5600[29])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i30_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i31_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [30]), 
         .D(key_mem_new[30]), .Z(key_mem_0__127__N_5600[30])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i31_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i32_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [31]), 
         .D(key_mem_new[31]), .Z(key_mem_0__127__N_5600[31])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i32_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i33_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [32]), 
         .D(key_mem_new[32]), .Z(key_mem_0__127__N_5600[32])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i33_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i34_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [33]), 
         .D(key_mem_new[33]), .Z(key_mem_0__127__N_5600[33])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i34_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i35_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [34]), 
         .D(key_mem_new[34]), .Z(key_mem_0__127__N_5600[34])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i35_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i36_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [35]), 
         .D(key_mem_new[35]), .Z(key_mem_0__127__N_5600[35])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i36_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i37_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [36]), 
         .D(key_mem_new[36]), .Z(key_mem_0__127__N_5600[36])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i37_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i38_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [37]), 
         .D(key_mem_new[37]), .Z(key_mem_0__127__N_5600[37])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i38_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i39_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [38]), 
         .D(key_mem_new[38]), .Z(key_mem_0__127__N_5600[38])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i39_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i40_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [39]), 
         .D(key_mem_new[39]), .Z(key_mem_0__127__N_5600[39])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i40_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i41_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [40]), 
         .D(key_mem_new[40]), .Z(key_mem_0__127__N_5600[40])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i41_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i42_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [41]), 
         .D(key_mem_new[41]), .Z(key_mem_0__127__N_5600[41])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i42_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i43_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [42]), 
         .D(key_mem_new[42]), .Z(key_mem_0__127__N_5600[42])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i43_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i44_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [43]), 
         .D(key_mem_new[43]), .Z(key_mem_0__127__N_5600[43])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i44_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i45_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [44]), 
         .D(key_mem_new[44]), .Z(key_mem_0__127__N_5600[44])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i45_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i46_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [45]), 
         .D(key_mem_new[45]), .Z(key_mem_0__127__N_5600[45])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i46_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i47_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [46]), 
         .D(key_mem_new[46]), .Z(key_mem_0__127__N_5600[46])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i47_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i48_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [47]), 
         .D(key_mem_new[47]), .Z(key_mem_0__127__N_5600[47])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i48_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i49_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [48]), 
         .D(key_mem_new[48]), .Z(key_mem_0__127__N_5600[48])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i49_3_lut_4_lut.init = 16'hf1e0;
    L6MUX21 i25879 (.D0(n31034), .D1(n31035), .SD(\muxed_round_nr[2] ), 
            .Z(n31038));
    L6MUX21 i25880 (.D0(n31036), .D1(n33384), .SD(\muxed_round_nr[2] ), 
            .Z(n31039));
    LUT4 i2_2_lut_rep_341 (.A(prev_key0_reg[75]), .B(n4_adj_8361), .Z(n33645)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i2_2_lut_rep_341.init = 16'h6666;
    L6MUX21 i25886 (.D0(n31041), .D1(n31042), .SD(\muxed_round_nr[2] ), 
            .Z(n31045));
    L6MUX21 i25887 (.D0(n31043), .D1(n33386), .SD(\muxed_round_nr[2] ), 
            .Z(n31046));
    LUT4 round_3__I_0_Mux_101_i11_3_lut (.A(\key_mem[12] [101]), .B(\key_mem[13] [101]), 
         .C(n33952), .Z(n11_adj_125)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_101_i11_3_lut.init = 16'hcaca;
    LUT4 mux_51_i108_3_lut_4_lut (.A(prev_key1_reg[107]), .B(\round_key_gen.trw[11] ), 
         .C(n33860), .D(\key_reg[0] [11]), .Z(key_mem_new_127__N_7264[107])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam mux_51_i108_3_lut_4_lut.init = 16'h6f60;
    L6MUX21 i25893 (.D0(n31048), .D1(n31049), .SD(\muxed_round_nr[2] ), 
            .Z(n31052));
    L6MUX21 i25894 (.D0(n31050), .D1(n33387), .SD(\muxed_round_nr[2] ), 
            .Z(n31053));
    L6MUX21 i25900 (.D0(n31055), .D1(n31056), .SD(\muxed_round_nr[2] ), 
            .Z(n31059));
    L6MUX21 i25901 (.D0(n31057), .D1(n33389), .SD(\muxed_round_nr[2] ), 
            .Z(n31060));
    LUT4 i3310_3_lut_4_lut (.A(prev_key1_reg[106]), .B(\round_key_gen.trw[10] ), 
         .C(n35835), .D(n33604), .Z(n8795)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam i3310_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_51_i107_3_lut_4_lut (.A(prev_key1_reg[106]), .B(\round_key_gen.trw[10] ), 
         .C(n33860), .D(\key_reg[0] [10]), .Z(key_mem_new_127__N_7264[106])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam mux_51_i107_3_lut_4_lut.init = 16'h6f60;
    L6MUX21 i25907 (.D0(n31062), .D1(n31063), .SD(\muxed_round_nr[2] ), 
            .Z(n31066));
    L6MUX21 i25908 (.D0(n31064), .D1(n33391), .SD(\muxed_round_nr[2] ), 
            .Z(n31067));
    L6MUX21 i25914 (.D0(n31069), .D1(n31070), .SD(\muxed_round_nr[2] ), 
            .Z(n31073));
    L6MUX21 i25915 (.D0(n31071), .D1(n33393), .SD(\muxed_round_nr[2] ), 
            .Z(n31074));
    LUT4 i3308_3_lut_4_lut (.A(prev_key1_reg[105]), .B(\round_key_gen.trw[9] ), 
         .C(n35835), .D(n33605), .Z(n8793)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam i3308_3_lut_4_lut.init = 16'hf606;
    L6MUX21 i25921 (.D0(n31076), .D1(n31077), .SD(\muxed_round_nr[2] ), 
            .Z(n31080));
    L6MUX21 i25922 (.D0(n31078), .D1(n33395), .SD(\muxed_round_nr[2] ), 
            .Z(n31081));
    L6MUX21 i25928 (.D0(n31083), .D1(n31084), .SD(\muxed_round_nr[2] ), 
            .Z(n31087));
    L6MUX21 i25929 (.D0(n31085), .D1(n33398), .SD(\muxed_round_nr[2] ), 
            .Z(n31088));
    LUT4 mux_51_i106_3_lut_4_lut (.A(prev_key1_reg[105]), .B(\round_key_gen.trw[9] ), 
         .C(n33860), .D(\key_reg[0] [9]), .Z(key_mem_new_127__N_7264[105])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam mux_51_i106_3_lut_4_lut.init = 16'h6f60;
    L6MUX21 i25935 (.D0(n31090), .D1(n31091), .SD(\muxed_round_nr[2] ), 
            .Z(n31094));
    L6MUX21 i25936 (.D0(n31092), .D1(n33400), .SD(\muxed_round_nr[2] ), 
            .Z(n31095));
    LUT4 round_3__I_0_Mux_101_i9_3_lut (.A(\key_mem[10] [101]), .B(\key_mem[11] [101]), 
         .C(n33952), .Z(n9_adj_9276)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_101_i9_3_lut.init = 16'hcaca;
    L6MUX21 i25942 (.D0(n31097), .D1(n31098), .SD(\muxed_round_nr[2] ), 
            .Z(n31101));
    L6MUX21 i25943 (.D0(n31099), .D1(n33402), .SD(\muxed_round_nr[2] ), 
            .Z(n31102));
    LUT4 round_3__I_0_Mux_101_i8_3_lut (.A(\key_mem[8] [101]), .B(\key_mem[9] [101]), 
         .C(n33952), .Z(n8_adj_9277)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_101_i8_3_lut.init = 16'hcaca;
    L6MUX21 i25949 (.D0(n31104), .D1(n31105), .SD(\muxed_round_nr[2] ), 
            .Z(n31108));
    L6MUX21 i25950 (.D0(n31106), .D1(n33405), .SD(\muxed_round_nr[2] ), 
            .Z(n31109));
    L6MUX21 i25956 (.D0(n31111), .D1(n31112), .SD(\muxed_round_nr[2] ), 
            .Z(n31115));
    L6MUX21 i25957 (.D0(n31113), .D1(n33406), .SD(\muxed_round_nr[2] ), 
            .Z(n31116));
    LUT4 i3306_3_lut_4_lut (.A(prev_key1_reg[104]), .B(\round_key_gen.trw[8] ), 
         .C(n35835), .D(n33606), .Z(n8791)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam i3306_3_lut_4_lut.init = 16'hf606;
    L6MUX21 i25963 (.D0(n31118), .D1(n31119), .SD(\muxed_round_nr[2] ), 
            .Z(n31122));
    L6MUX21 i25964 (.D0(n31120), .D1(n33409), .SD(\muxed_round_nr[2] ), 
            .Z(n31123));
    LUT4 round_3__I_0_Mux_101_i5_3_lut (.A(\key_mem[6] [101]), .B(\key_mem[7] [101]), 
         .C(n33952), .Z(n5_adj_9278)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_101_i5_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_101_i4_3_lut (.A(\key_mem[4] [101]), .B(\key_mem[5] [101]), 
         .C(n33952), .Z(n4_adj_9279)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_101_i4_3_lut.init = 16'hcaca;
    L6MUX21 i25970 (.D0(n31125), .D1(n31126), .SD(\muxed_round_nr[2] ), 
            .Z(n31129));
    L6MUX21 i25971 (.D0(n31127), .D1(n33411), .SD(\muxed_round_nr[2] ), 
            .Z(n31130));
    LUT4 mux_51_i105_3_lut_4_lut (.A(prev_key1_reg[104]), .B(\round_key_gen.trw[8] ), 
         .C(n33860), .D(\key_reg[0] [8]), .Z(key_mem_new_127__N_7264[104])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam mux_51_i105_3_lut_4_lut.init = 16'h6f60;
    LUT4 i3304_3_lut_4_lut (.A(prev_key1_reg[103]), .B(\round_key_gen.trw[7] ), 
         .C(n35835), .D(n33607), .Z(n8789)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam i3304_3_lut_4_lut.init = 16'hf606;
    L6MUX21 i25977 (.D0(n31132), .D1(n31133), .SD(\muxed_round_nr[2] ), 
            .Z(n31136));
    L6MUX21 i25978 (.D0(n31134), .D1(n33413), .SD(\muxed_round_nr[2] ), 
            .Z(n31137));
    LUT4 mux_51_i104_3_lut_4_lut (.A(prev_key1_reg[103]), .B(\round_key_gen.trw[7] ), 
         .C(n33860), .D(\key_reg[0] [7]), .Z(key_mem_new_127__N_7264[103])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam mux_51_i104_3_lut_4_lut.init = 16'h6f60;
    PFUMX i25861 (.BLUT(n1_adj_9214), .ALUT(n2_adj_9213), .C0(\muxed_round_nr[1] ), 
          .Z(n31020));
    LUT4 round_3__I_0_Mux_101_i2_3_lut (.A(\key_mem[2] [101]), .B(\key_mem[3] [101]), 
         .C(n33952), .Z(n2_adj_9280)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_101_i2_3_lut.init = 16'hcaca;
    PFUMX i24988 (.BLUT(n1_adj_9212), .ALUT(n2_adj_9211), .C0(\muxed_round_nr[1] ), 
          .Z(n30147));
    LUT4 i3302_3_lut_4_lut (.A(prev_key1_reg[102]), .B(\round_key_gen.trw[6] ), 
         .C(n35835), .D(n33608), .Z(n8787)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam i3302_3_lut_4_lut.init = 16'hf606;
    LUT4 round_3__I_0_Mux_101_i1_3_lut (.A(\key_mem[0] [101]), .B(\key_mem[1] [101]), 
         .C(n33952), .Z(n1_adj_9281)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_101_i1_3_lut.init = 16'hcaca;
    PFUMX i24989 (.BLUT(n4_adj_9210), .ALUT(n5_adj_9209), .C0(\muxed_round_nr[1] ), 
          .Z(n30148));
    LUT4 mux_51_i103_3_lut_4_lut (.A(prev_key1_reg[102]), .B(\round_key_gen.trw[6] ), 
         .C(n33860), .D(\key_reg[0] [6]), .Z(key_mem_new_127__N_7264[102])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam mux_51_i103_3_lut_4_lut.init = 16'h6f60;
    PFUMX i24990 (.BLUT(n8_adj_9208), .ALUT(n9_adj_9207), .C0(\muxed_round_nr[1] ), 
          .Z(n30149));
    LUT4 i3300_3_lut_4_lut (.A(prev_key1_reg[101]), .B(\round_key_gen.trw[5] ), 
         .C(n35835), .D(n33609), .Z(n8785)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam i3300_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_85_i76_3_lut_rep_242_4_lut (.A(prev_key0_reg[75]), .B(n4_adj_8361), 
         .C(n33859), .D(\key_reg[5] [11]), .Z(n33546)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam mux_85_i76_3_lut_rep_242_4_lut.init = 16'h6f60;
    LUT4 mux_51_i102_3_lut_4_lut (.A(prev_key1_reg[101]), .B(\round_key_gen.trw[5] ), 
         .C(n33860), .D(\key_reg[0] [5]), .Z(key_mem_new_127__N_7264[101])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam mux_51_i102_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_18_i50_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [49]), 
         .D(key_mem_new[49]), .Z(key_mem_0__127__N_5600[49])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i50_3_lut_4_lut.init = 16'hf1e0;
    LUT4 round_3__I_0_Mux_100_i11_3_lut (.A(\key_mem[12] [100]), .B(\key_mem[13] [100]), 
         .C(n33952), .Z(n11_adj_126)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_100_i11_3_lut.init = 16'hcaca;
    LUT4 mux_18_i51_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [50]), 
         .D(key_mem_new[50]), .Z(key_mem_0__127__N_5600[50])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i51_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i24995 (.BLUT(n1_adj_9204), .ALUT(n2_adj_9203), .C0(\muxed_round_nr[1] ), 
          .Z(n30154));
    PFUMX i25718 (.BLUT(n8_adj_9205), .ALUT(n9_adj_9163), .C0(\muxed_round_nr[1] ), 
          .Z(n30877));
    LUT4 mux_18_i52_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [51]), 
         .D(key_mem_new[51]), .Z(key_mem_0__127__N_5600[51])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i52_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i53_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [52]), 
         .D(key_mem_new[52]), .Z(key_mem_0__127__N_5600[52])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i53_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3298_3_lut_4_lut (.A(prev_key1_reg[100]), .B(\round_key_gen.trw[4] ), 
         .C(n35835), .D(n33610), .Z(n8783)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam i3298_3_lut_4_lut.init = 16'hf606;
    PFUMX i24996 (.BLUT(n4_adj_9202), .ALUT(n5_adj_9201), .C0(\muxed_round_nr[1] ), 
          .Z(n30155));
    PFUMX i24997 (.BLUT(n8_adj_9200), .ALUT(n9_adj_9199), .C0(\muxed_round_nr[1] ), 
          .Z(n30156));
    LUT4 round_3__I_0_Mux_100_i9_3_lut (.A(\key_mem[10] [100]), .B(\key_mem[11] [100]), 
         .C(n33952), .Z(n9_adj_9283)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_100_i9_3_lut.init = 16'hcaca;
    LUT4 mux_18_i54_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [53]), 
         .D(key_mem_new[53]), .Z(key_mem_0__127__N_5600[53])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i54_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25002 (.BLUT(n1_adj_9197), .ALUT(n2_adj_9196), .C0(\muxed_round_nr[1] ), 
          .Z(n30161));
    LUT4 mux_18_i55_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [54]), 
         .D(key_mem_new[54]), .Z(key_mem_0__127__N_5600[54])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i55_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_51_i101_3_lut_4_lut (.A(prev_key1_reg[100]), .B(\round_key_gen.trw[4] ), 
         .C(n33860), .D(\key_reg[0] [4]), .Z(key_mem_new_127__N_7264[100])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam mux_51_i101_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_18_i56_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [55]), 
         .D(key_mem_new[55]), .Z(key_mem_0__127__N_5600[55])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i56_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25003 (.BLUT(n4_adj_9195), .ALUT(n5_adj_9194), .C0(\muxed_round_nr[1] ), 
          .Z(n30162));
    LUT4 round_3__I_0_Mux_100_i8_3_lut (.A(\key_mem[8] [100]), .B(\key_mem[9] [100]), 
         .C(n33952), .Z(n8_adj_9284)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_100_i8_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_100_i5_3_lut (.A(\key_mem[6] [100]), .B(\key_mem[7] [100]), 
         .C(n33952), .Z(n5_adj_9285)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_100_i5_3_lut.init = 16'hcaca;
    PFUMX i25004 (.BLUT(n8_adj_9193), .ALUT(n9_adj_9192), .C0(\muxed_round_nr[1] ), 
          .Z(n30163));
    LUT4 i3296_3_lut_4_lut (.A(prev_key1_reg[99]), .B(\round_key_gen.trw[3] ), 
         .C(n35835), .D(n33611), .Z(n8781)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam i3296_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_18_i57_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [56]), 
         .D(key_mem_new[56]), .Z(key_mem_0__127__N_5600[56])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i57_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i6_2_lut_3_lut_adj_663 (.A(prev_key1_reg[42]), .B(n33737), .C(keymem_sboxw[10]), 
         .Z(n15957)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;
    defparam i6_2_lut_3_lut_adj_663.init = 16'h9696;
    PFUMX i25009 (.BLUT(n1_adj_9190), .ALUT(n2_adj_9189), .C0(\muxed_round_nr[1] ), 
          .Z(n30168));
    PFUMX i25010 (.BLUT(n4_adj_9188), .ALUT(n5_adj_9187), .C0(\muxed_round_nr[1] ), 
          .Z(n30169));
    LUT4 mux_51_i100_3_lut_4_lut (.A(prev_key1_reg[99]), .B(\round_key_gen.trw[3] ), 
         .C(n33860), .D(\key_reg[0] [3]), .Z(key_mem_new_127__N_7264[99])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam mux_51_i100_3_lut_4_lut.init = 16'h6f60;
    LUT4 round_3__I_0_Mux_100_i4_3_lut (.A(\key_mem[4] [100]), .B(\key_mem[5] [100]), 
         .C(n33952), .Z(n4_adj_9286)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_100_i4_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_100_i2_3_lut (.A(\key_mem[2] [100]), .B(\key_mem[3] [100]), 
         .C(n33952), .Z(n2_adj_9287)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_100_i2_3_lut.init = 16'hcaca;
    PFUMX i25011 (.BLUT(n8_adj_9186), .ALUT(n9_adj_9185), .C0(\muxed_round_nr[1] ), 
          .Z(n30170));
    LUT4 i3294_3_lut_4_lut (.A(prev_key1_reg[98]), .B(\round_key_gen.trw[2] ), 
         .C(n35835), .D(n33612), .Z(n8779)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(244[26:34])
    defparam i3294_3_lut_4_lut.init = 16'hf606;
    PFUMX i25016 (.BLUT(n1_adj_9183), .ALUT(n2_adj_9182), .C0(\muxed_round_nr[1] ), 
          .Z(n30175));
    LUT4 round_3__I_0_Mux_100_i1_3_lut (.A(\key_mem[0] [100]), .B(\key_mem[1] [100]), 
         .C(n33952), .Z(n1_adj_9288)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_100_i1_3_lut.init = 16'hcaca;
    PFUMX i25017 (.BLUT(n4_adj_9181), .ALUT(n5_adj_9180), .C0(\muxed_round_nr[1] ), 
          .Z(n30176));
    LUT4 mux_18_i58_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [57]), 
         .D(key_mem_new[57]), .Z(key_mem_0__127__N_5600[57])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i58_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i59_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [58]), 
         .D(key_mem_new[58]), .Z(key_mem_0__127__N_5600[58])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i59_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i60_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [59]), 
         .D(key_mem_new[59]), .Z(key_mem_0__127__N_5600[59])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i60_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i61_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [60]), 
         .D(key_mem_new[60]), .Z(key_mem_0__127__N_5600[60])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i61_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25018 (.BLUT(n8_adj_9179), .ALUT(n9_adj_9178), .C0(\muxed_round_nr[1] ), 
          .Z(n30177));
    LUT4 mux_18_i62_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [61]), 
         .D(key_mem_new[61]), .Z(key_mem_0__127__N_5600[61])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i62_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i63_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [62]), 
         .D(key_mem_new[62]), .Z(key_mem_0__127__N_5600[62])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i63_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i64_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [63]), 
         .D(key_mem_new[63]), .Z(key_mem_0__127__N_5600[63])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i64_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i65_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [64]), 
         .D(key_mem_new[64]), .Z(key_mem_0__127__N_5600[64])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i65_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i66_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [65]), 
         .D(key_mem_new[65]), .Z(key_mem_0__127__N_5600[65])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i66_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i67_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [66]), 
         .D(key_mem_new[66]), .Z(key_mem_0__127__N_5600[66])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i67_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25023 (.BLUT(n1_adj_9176), .ALUT(n2_adj_9175), .C0(\muxed_round_nr[1] ), 
          .Z(n30182));
    LUT4 mux_18_i68_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [67]), 
         .D(key_mem_new[67]), .Z(key_mem_0__127__N_5600[67])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i68_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i69_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [68]), 
         .D(key_mem_new[68]), .Z(key_mem_0__127__N_5600[68])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i69_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25024 (.BLUT(n4_adj_9174), .ALUT(n5_adj_9173), .C0(\muxed_round_nr[1] ), 
          .Z(n30183));
    LUT4 mux_18_i70_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [69]), 
         .D(key_mem_new[69]), .Z(key_mem_0__127__N_5600[69])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i70_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i71_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [70]), 
         .D(key_mem_new[70]), .Z(key_mem_0__127__N_5600[70])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i71_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i72_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [71]), 
         .D(key_mem_new[71]), .Z(key_mem_0__127__N_5600[71])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i72_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i73_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [72]), 
         .D(key_mem_new[72]), .Z(key_mem_0__127__N_5600[72])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i73_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25025 (.BLUT(n8_adj_9172), .ALUT(n9_adj_9171), .C0(\muxed_round_nr[1] ), 
          .Z(n30184));
    LUT4 mux_18_i74_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [73]), 
         .D(key_mem_new[73]), .Z(key_mem_0__127__N_5600[73])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i74_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i75_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [74]), 
         .D(key_mem_new[74]), .Z(key_mem_0__127__N_5600[74])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i75_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i76_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [75]), 
         .D(key_mem_new[75]), .Z(key_mem_0__127__N_5600[75])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i76_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i77_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [76]), 
         .D(key_mem_new[76]), .Z(key_mem_0__127__N_5600[76])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i77_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25030 (.BLUT(n1_adj_9169), .ALUT(n2_adj_9168), .C0(\muxed_round_nr[1] ), 
          .Z(n30189));
    LUT4 mux_18_i78_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [77]), 
         .D(key_mem_new[77]), .Z(key_mem_0__127__N_5600[77])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i78_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25031 (.BLUT(n4_adj_9167), .ALUT(n5_adj_9166), .C0(\muxed_round_nr[1] ), 
          .Z(n30190));
    LUT4 mux_18_i79_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [78]), 
         .D(key_mem_new[78]), .Z(key_mem_0__127__N_5600[78])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i79_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i80_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [79]), 
         .D(key_mem_new[79]), .Z(key_mem_0__127__N_5600[79])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i80_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i81_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [80]), 
         .D(key_mem_new[80]), .Z(key_mem_0__127__N_5600[80])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i81_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25032 (.BLUT(n8_adj_9165), .ALUT(n9_adj_9164), .C0(\muxed_round_nr[1] ), 
          .Z(n30191));
    LUT4 mux_18_i82_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [81]), 
         .D(key_mem_new[81]), .Z(key_mem_0__127__N_5600[81])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i82_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i83_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [82]), 
         .D(key_mem_new[82]), .Z(key_mem_0__127__N_5600[82])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i83_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i84_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [83]), 
         .D(key_mem_new[83]), .Z(key_mem_0__127__N_5600[83])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i84_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i85_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [84]), 
         .D(key_mem_new[84]), .Z(key_mem_0__127__N_5600[84])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i85_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i86_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [85]), 
         .D(key_mem_new[85]), .Z(key_mem_0__127__N_5600[85])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i86_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i87_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [86]), 
         .D(key_mem_new[86]), .Z(key_mem_0__127__N_5600[86])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i87_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i88_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [87]), 
         .D(key_mem_new[87]), .Z(key_mem_0__127__N_5600[87])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i88_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i89_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [88]), 
         .D(key_mem_new[88]), .Z(key_mem_0__127__N_5600[88])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i89_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i90_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [89]), 
         .D(key_mem_new[89]), .Z(key_mem_0__127__N_5600[89])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i90_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i91_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [90]), 
         .D(key_mem_new[90]), .Z(key_mem_0__127__N_5600[90])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i91_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i92_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [91]), 
         .D(key_mem_new[91]), .Z(key_mem_0__127__N_5600[91])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i92_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i93_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [92]), 
         .D(key_mem_new[92]), .Z(key_mem_0__127__N_5600[92])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i93_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i94_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [93]), 
         .D(key_mem_new[93]), .Z(key_mem_0__127__N_5600[93])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i94_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i95_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [94]), 
         .D(key_mem_new[94]), .Z(key_mem_0__127__N_5600[94])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i95_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i96_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [95]), 
         .D(key_mem_new[95]), .Z(key_mem_0__127__N_5600[95])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i96_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i97_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [96]), 
         .D(key_mem_new[96]), .Z(key_mem_0__127__N_5600[96])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i97_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i98_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [97]), 
         .D(key_mem_new[97]), .Z(key_mem_0__127__N_5600[97])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i98_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i99_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [98]), 
         .D(key_mem_new[98]), .Z(key_mem_0__127__N_5600[98])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i99_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i100_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [99]), 
         .D(key_mem_new[99]), .Z(key_mem_0__127__N_5600[99])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i100_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i101_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [100]), 
         .D(key_mem_new[100]), .Z(key_mem_0__127__N_5600[100])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i101_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i102_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [101]), 
         .D(key_mem_new[101]), .Z(key_mem_0__127__N_5600[101])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i102_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i103_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [102]), 
         .D(key_mem_new[102]), .Z(key_mem_0__127__N_5600[102])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i103_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i104_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [103]), 
         .D(key_mem_new[103]), .Z(key_mem_0__127__N_5600[103])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i104_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i105_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [104]), 
         .D(key_mem_new[104]), .Z(key_mem_0__127__N_5600[104])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i105_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i106_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [105]), 
         .D(key_mem_new[105]), .Z(key_mem_0__127__N_5600[105])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i106_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i107_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [106]), 
         .D(key_mem_new[106]), .Z(key_mem_0__127__N_5600[106])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i107_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i108_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [107]), 
         .D(key_mem_new[107]), .Z(key_mem_0__127__N_5600[107])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i108_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i109_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [108]), 
         .D(key_mem_new[108]), .Z(key_mem_0__127__N_5600[108])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i109_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i110_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [109]), 
         .D(key_mem_new[109]), .Z(key_mem_0__127__N_5600[109])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i110_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i111_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [110]), 
         .D(key_mem_new[110]), .Z(key_mem_0__127__N_5600[110])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i111_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i112_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [111]), 
         .D(key_mem_new[111]), .Z(key_mem_0__127__N_5600[111])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i112_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i113_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [112]), 
         .D(key_mem_new[112]), .Z(key_mem_0__127__N_5600[112])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i113_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i114_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [113]), 
         .D(key_mem_new[113]), .Z(key_mem_0__127__N_5600[113])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i114_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i115_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [114]), 
         .D(key_mem_new[114]), .Z(key_mem_0__127__N_5600[114])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i115_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i116_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [115]), 
         .D(key_mem_new[115]), .Z(key_mem_0__127__N_5600[115])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i116_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i117_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [116]), 
         .D(key_mem_new[116]), .Z(key_mem_0__127__N_5600[116])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i117_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i118_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [117]), 
         .D(key_mem_new[117]), .Z(key_mem_0__127__N_5600[117])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i118_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i119_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [118]), 
         .D(key_mem_new[118]), .Z(key_mem_0__127__N_5600[118])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i119_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i120_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [119]), 
         .D(key_mem_new[119]), .Z(key_mem_0__127__N_5600[119])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i120_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i121_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [120]), 
         .D(key_mem_new[120]), .Z(key_mem_0__127__N_5600[120])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i121_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i122_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [121]), 
         .D(key_mem_new[121]), .Z(key_mem_0__127__N_5600[121])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i122_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i123_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [122]), 
         .D(key_mem_new[122]), .Z(key_mem_0__127__N_5600[122])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i123_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i124_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [123]), 
         .D(key_mem_new[123]), .Z(key_mem_0__127__N_5600[123])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i124_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i125_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [124]), 
         .D(key_mem_new[124]), .Z(key_mem_0__127__N_5600[124])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i125_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i126_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [125]), 
         .D(key_mem_new[125]), .Z(key_mem_0__127__N_5600[125])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i126_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i127_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [126]), 
         .D(key_mem_new[126]), .Z(key_mem_0__127__N_5600[126])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i127_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_18_i128_3_lut_4_lut (.A(n33945), .B(n33916), .C(\key_mem[5] [127]), 
         .D(key_mem_new[127]), .Z(key_mem_0__127__N_5600[127])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_18_i128_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i1_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [0]), 
         .D(key_mem_new[0]), .Z(key_mem_0__127__N_5728[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i2_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [1]), 
         .D(key_mem_new[1]), .Z(key_mem_0__127__N_5728[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i3_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [2]), 
         .D(key_mem_new[2]), .Z(key_mem_0__127__N_5728[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i4_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [3]), 
         .D(key_mem_new[3]), .Z(key_mem_0__127__N_5728[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i5_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [4]), 
         .D(key_mem_new[4]), .Z(key_mem_0__127__N_5728[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i6_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [5]), 
         .D(key_mem_new[5]), .Z(key_mem_0__127__N_5728[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i7_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [6]), 
         .D(key_mem_new[6]), .Z(key_mem_0__127__N_5728[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i8_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [7]), 
         .D(key_mem_new[7]), .Z(key_mem_0__127__N_5728[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i9_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [8]), 
         .D(key_mem_new[8]), .Z(key_mem_0__127__N_5728[8])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i9_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i10_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [9]), 
         .D(key_mem_new[9]), .Z(key_mem_0__127__N_5728[9])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i10_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i11_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [10]), 
         .D(key_mem_new[10]), .Z(key_mem_0__127__N_5728[10])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i11_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i12_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [11]), 
         .D(key_mem_new[11]), .Z(key_mem_0__127__N_5728[11])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i12_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i13_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [12]), 
         .D(key_mem_new[12]), .Z(key_mem_0__127__N_5728[12])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i13_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i14_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [13]), 
         .D(key_mem_new[13]), .Z(key_mem_0__127__N_5728[13])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i14_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i15_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [14]), 
         .D(key_mem_new[14]), .Z(key_mem_0__127__N_5728[14])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i15_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i16_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [15]), 
         .D(key_mem_new[15]), .Z(key_mem_0__127__N_5728[15])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i16_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i17_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [16]), 
         .D(key_mem_new[16]), .Z(key_mem_0__127__N_5728[16])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i17_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i18_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [17]), 
         .D(key_mem_new[17]), .Z(key_mem_0__127__N_5728[17])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i18_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i19_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [18]), 
         .D(key_mem_new[18]), .Z(key_mem_0__127__N_5728[18])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i19_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i20_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [19]), 
         .D(key_mem_new[19]), .Z(key_mem_0__127__N_5728[19])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i20_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i21_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [20]), 
         .D(key_mem_new[20]), .Z(key_mem_0__127__N_5728[20])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i21_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i22_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [21]), 
         .D(key_mem_new[21]), .Z(key_mem_0__127__N_5728[21])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i22_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i23_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [22]), 
         .D(key_mem_new[22]), .Z(key_mem_0__127__N_5728[22])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i23_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i24_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [23]), 
         .D(key_mem_new[23]), .Z(key_mem_0__127__N_5728[23])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i24_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i25_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [24]), 
         .D(key_mem_new[24]), .Z(key_mem_0__127__N_5728[24])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i25_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i26_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [25]), 
         .D(key_mem_new[25]), .Z(key_mem_0__127__N_5728[25])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i26_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i27_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [26]), 
         .D(key_mem_new[26]), .Z(key_mem_0__127__N_5728[26])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i27_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i28_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [27]), 
         .D(key_mem_new[27]), .Z(key_mem_0__127__N_5728[27])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i28_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i29_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [28]), 
         .D(key_mem_new[28]), .Z(key_mem_0__127__N_5728[28])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i29_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i30_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [29]), 
         .D(key_mem_new[29]), .Z(key_mem_0__127__N_5728[29])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i30_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i31_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [30]), 
         .D(key_mem_new[30]), .Z(key_mem_0__127__N_5728[30])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i31_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i32_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [31]), 
         .D(key_mem_new[31]), .Z(key_mem_0__127__N_5728[31])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i32_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i33_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [32]), 
         .D(key_mem_new[32]), .Z(key_mem_0__127__N_5728[32])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i33_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i34_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [33]), 
         .D(key_mem_new[33]), .Z(key_mem_0__127__N_5728[33])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i34_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i35_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [34]), 
         .D(key_mem_new[34]), .Z(key_mem_0__127__N_5728[34])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i35_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i36_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [35]), 
         .D(key_mem_new[35]), .Z(key_mem_0__127__N_5728[35])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i36_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i37_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [36]), 
         .D(key_mem_new[36]), .Z(key_mem_0__127__N_5728[36])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i37_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i38_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [37]), 
         .D(key_mem_new[37]), .Z(key_mem_0__127__N_5728[37])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i38_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i39_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [38]), 
         .D(key_mem_new[38]), .Z(key_mem_0__127__N_5728[38])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i39_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i40_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [39]), 
         .D(key_mem_new[39]), .Z(key_mem_0__127__N_5728[39])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i40_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i41_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [40]), 
         .D(key_mem_new[40]), .Z(key_mem_0__127__N_5728[40])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i41_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i42_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [41]), 
         .D(key_mem_new[41]), .Z(key_mem_0__127__N_5728[41])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i42_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i43_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [42]), 
         .D(key_mem_new[42]), .Z(key_mem_0__127__N_5728[42])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i43_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i44_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [43]), 
         .D(key_mem_new[43]), .Z(key_mem_0__127__N_5728[43])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i44_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i45_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [44]), 
         .D(key_mem_new[44]), .Z(key_mem_0__127__N_5728[44])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i45_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i46_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [45]), 
         .D(key_mem_new[45]), .Z(key_mem_0__127__N_5728[45])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i46_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i47_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [46]), 
         .D(key_mem_new[46]), .Z(key_mem_0__127__N_5728[46])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i47_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i48_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [47]), 
         .D(key_mem_new[47]), .Z(key_mem_0__127__N_5728[47])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i48_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i49_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [48]), 
         .D(key_mem_new[48]), .Z(key_mem_0__127__N_5728[48])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i49_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i50_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [49]), 
         .D(key_mem_new[49]), .Z(key_mem_0__127__N_5728[49])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i50_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i51_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [50]), 
         .D(key_mem_new[50]), .Z(key_mem_0__127__N_5728[50])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i51_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i52_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [51]), 
         .D(key_mem_new[51]), .Z(key_mem_0__127__N_5728[51])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i52_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i53_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [52]), 
         .D(key_mem_new[52]), .Z(key_mem_0__127__N_5728[52])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i53_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i54_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [53]), 
         .D(key_mem_new[53]), .Z(key_mem_0__127__N_5728[53])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i54_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i55_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [54]), 
         .D(key_mem_new[54]), .Z(key_mem_0__127__N_5728[54])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i55_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i56_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [55]), 
         .D(key_mem_new[55]), .Z(key_mem_0__127__N_5728[55])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i56_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i57_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [56]), 
         .D(key_mem_new[56]), .Z(key_mem_0__127__N_5728[56])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i57_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i58_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [57]), 
         .D(key_mem_new[57]), .Z(key_mem_0__127__N_5728[57])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i58_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i59_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [58]), 
         .D(key_mem_new[58]), .Z(key_mem_0__127__N_5728[58])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i59_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i60_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [59]), 
         .D(key_mem_new[59]), .Z(key_mem_0__127__N_5728[59])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i60_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i61_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [60]), 
         .D(key_mem_new[60]), .Z(key_mem_0__127__N_5728[60])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i61_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i62_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [61]), 
         .D(key_mem_new[61]), .Z(key_mem_0__127__N_5728[61])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i62_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i63_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [62]), 
         .D(key_mem_new[62]), .Z(key_mem_0__127__N_5728[62])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i63_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i64_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [63]), 
         .D(key_mem_new[63]), .Z(key_mem_0__127__N_5728[63])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i64_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i65_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [64]), 
         .D(key_mem_new[64]), .Z(key_mem_0__127__N_5728[64])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i65_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i66_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [65]), 
         .D(key_mem_new[65]), .Z(key_mem_0__127__N_5728[65])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i66_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i67_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [66]), 
         .D(key_mem_new[66]), .Z(key_mem_0__127__N_5728[66])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i67_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i68_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [67]), 
         .D(key_mem_new[67]), .Z(key_mem_0__127__N_5728[67])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i68_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i69_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [68]), 
         .D(key_mem_new[68]), .Z(key_mem_0__127__N_5728[68])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i69_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i70_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [69]), 
         .D(key_mem_new[69]), .Z(key_mem_0__127__N_5728[69])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i70_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i71_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [70]), 
         .D(key_mem_new[70]), .Z(key_mem_0__127__N_5728[70])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i71_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i72_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [71]), 
         .D(key_mem_new[71]), .Z(key_mem_0__127__N_5728[71])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i72_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i73_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [72]), 
         .D(key_mem_new[72]), .Z(key_mem_0__127__N_5728[72])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i73_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i74_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [73]), 
         .D(key_mem_new[73]), .Z(key_mem_0__127__N_5728[73])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i74_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i75_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [74]), 
         .D(key_mem_new[74]), .Z(key_mem_0__127__N_5728[74])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i75_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i76_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [75]), 
         .D(key_mem_new[75]), .Z(key_mem_0__127__N_5728[75])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i76_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i77_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [76]), 
         .D(key_mem_new[76]), .Z(key_mem_0__127__N_5728[76])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i77_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i78_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [77]), 
         .D(key_mem_new[77]), .Z(key_mem_0__127__N_5728[77])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i78_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i79_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [78]), 
         .D(key_mem_new[78]), .Z(key_mem_0__127__N_5728[78])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i79_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i80_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [79]), 
         .D(key_mem_new[79]), .Z(key_mem_0__127__N_5728[79])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i80_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i81_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [80]), 
         .D(key_mem_new[80]), .Z(key_mem_0__127__N_5728[80])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i81_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i82_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [81]), 
         .D(key_mem_new[81]), .Z(key_mem_0__127__N_5728[81])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i82_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i83_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [82]), 
         .D(key_mem_new[82]), .Z(key_mem_0__127__N_5728[82])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i83_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i84_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [83]), 
         .D(key_mem_new[83]), .Z(key_mem_0__127__N_5728[83])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i84_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i85_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [84]), 
         .D(key_mem_new[84]), .Z(key_mem_0__127__N_5728[84])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i85_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i86_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [85]), 
         .D(key_mem_new[85]), .Z(key_mem_0__127__N_5728[85])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i86_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i87_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [86]), 
         .D(key_mem_new[86]), .Z(key_mem_0__127__N_5728[86])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i87_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i88_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [87]), 
         .D(key_mem_new[87]), .Z(key_mem_0__127__N_5728[87])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i88_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i89_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [88]), 
         .D(key_mem_new[88]), .Z(key_mem_0__127__N_5728[88])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i89_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25037 (.BLUT(n1_adj_9161), .ALUT(n2_adj_9160), .C0(\muxed_round_nr[1] ), 
          .Z(n30196));
    LUT4 mux_17_i90_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [89]), 
         .D(key_mem_new[89]), .Z(key_mem_0__127__N_5728[89])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i90_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i91_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [90]), 
         .D(key_mem_new[90]), .Z(key_mem_0__127__N_5728[90])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i91_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25038 (.BLUT(n4_adj_9159), .ALUT(n5_adj_9158), .C0(\muxed_round_nr[1] ), 
          .Z(n30197));
    LUT4 mux_17_i92_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [91]), 
         .D(key_mem_new[91]), .Z(key_mem_0__127__N_5728[91])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i92_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i93_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [92]), 
         .D(key_mem_new[92]), .Z(key_mem_0__127__N_5728[92])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i93_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i94_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [93]), 
         .D(key_mem_new[93]), .Z(key_mem_0__127__N_5728[93])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i94_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25039 (.BLUT(n8_adj_9157), .ALUT(n9_adj_9156), .C0(\muxed_round_nr[1] ), 
          .Z(n30198));
    LUT4 mux_17_i95_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [94]), 
         .D(key_mem_new[94]), .Z(key_mem_0__127__N_5728[94])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i95_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i96_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [95]), 
         .D(key_mem_new[95]), .Z(key_mem_0__127__N_5728[95])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i96_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i97_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [96]), 
         .D(key_mem_new[96]), .Z(key_mem_0__127__N_5728[96])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i97_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i98_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [97]), 
         .D(key_mem_new[97]), .Z(key_mem_0__127__N_5728[97])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i98_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i99_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [98]), 
         .D(key_mem_new[98]), .Z(key_mem_0__127__N_5728[98])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i99_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i100_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [99]), 
         .D(key_mem_new[99]), .Z(key_mem_0__127__N_5728[99])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i100_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25723 (.BLUT(n1_adj_9151), .ALUT(n2_adj_9145), .C0(\muxed_round_nr[1] ), 
          .Z(n30882));
    LUT4 mux_17_i101_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [100]), 
         .D(key_mem_new[100]), .Z(key_mem_0__127__N_5728[100])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i101_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i102_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [101]), 
         .D(key_mem_new[101]), .Z(key_mem_0__127__N_5728[101])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i102_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25044 (.BLUT(n1_adj_9153), .ALUT(n2_adj_9152), .C0(\muxed_round_nr[1] ), 
          .Z(n30203));
    LUT4 mux_17_i103_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [102]), 
         .D(key_mem_new[102]), .Z(key_mem_0__127__N_5728[102])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i103_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i104_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [103]), 
         .D(key_mem_new[103]), .Z(key_mem_0__127__N_5728[103])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i104_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i105_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [104]), 
         .D(key_mem_new[104]), .Z(key_mem_0__127__N_5728[104])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i105_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25045 (.BLUT(n4_adj_9150), .ALUT(n5_adj_9149), .C0(\muxed_round_nr[1] ), 
          .Z(n30204));
    LUT4 mux_17_i106_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [105]), 
         .D(key_mem_new[105]), .Z(key_mem_0__127__N_5728[105])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i106_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25046 (.BLUT(n8_adj_9148), .ALUT(n9_adj_9147), .C0(\muxed_round_nr[1] ), 
          .Z(n30205));
    LUT4 mux_17_i107_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [106]), 
         .D(key_mem_new[106]), .Z(key_mem_0__127__N_5728[106])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i107_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i108_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [107]), 
         .D(key_mem_new[107]), .Z(key_mem_0__127__N_5728[107])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i108_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i109_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [108]), 
         .D(key_mem_new[108]), .Z(key_mem_0__127__N_5728[108])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i109_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i110_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [109]), 
         .D(key_mem_new[109]), .Z(key_mem_0__127__N_5728[109])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i110_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i111_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [110]), 
         .D(key_mem_new[110]), .Z(key_mem_0__127__N_5728[110])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i111_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i112_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [111]), 
         .D(key_mem_new[111]), .Z(key_mem_0__127__N_5728[111])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i112_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i113_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [112]), 
         .D(key_mem_new[112]), .Z(key_mem_0__127__N_5728[112])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i113_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i114_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [113]), 
         .D(key_mem_new[113]), .Z(key_mem_0__127__N_5728[113])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i114_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25051 (.BLUT(n1_adj_9144), .ALUT(n2_adj_9143), .C0(\muxed_round_nr[1] ), 
          .Z(n30210));
    LUT4 mux_17_i115_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [114]), 
         .D(key_mem_new[114]), .Z(key_mem_0__127__N_5728[114])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i115_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i116_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [115]), 
         .D(key_mem_new[115]), .Z(key_mem_0__127__N_5728[115])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i116_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i117_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [116]), 
         .D(key_mem_new[116]), .Z(key_mem_0__127__N_5728[116])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i117_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25724 (.BLUT(n4_adj_9137), .ALUT(n5_adj_9129), .C0(\muxed_round_nr[1] ), 
          .Z(n30883));
    LUT4 mux_17_i118_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [117]), 
         .D(key_mem_new[117]), .Z(key_mem_0__127__N_5728[117])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i118_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i119_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [118]), 
         .D(key_mem_new[118]), .Z(key_mem_0__127__N_5728[118])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i119_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25052 (.BLUT(n4_adj_9142), .ALUT(n5_adj_9141), .C0(\muxed_round_nr[1] ), 
          .Z(n30211));
    LUT4 mux_17_i120_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [119]), 
         .D(key_mem_new[119]), .Z(key_mem_0__127__N_5728[119])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i120_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25053 (.BLUT(n8_adj_9140), .ALUT(n9_adj_9139), .C0(\muxed_round_nr[1] ), 
          .Z(n30212));
    LUT4 mux_17_i121_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [120]), 
         .D(key_mem_new[120]), .Z(key_mem_0__127__N_5728[120])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i121_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i122_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [121]), 
         .D(key_mem_new[121]), .Z(key_mem_0__127__N_5728[121])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i122_3_lut_4_lut.init = 16'hf1e0;
    FD1P3IX round_ctr_reg_912__i3 (.D(n3[3]), .SP(round_ctr_we), .CD(n6361[2]), 
            .CK(clk_c), .Q(round_ctr_reg[3]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(352[27:47])
    defparam round_ctr_reg_912__i3.GSR = "ENABLED";
    FD1P3IX round_ctr_reg_912__i2 (.D(n3[2]), .SP(round_ctr_we), .CD(n6361[2]), 
            .CK(clk_c), .Q(round_ctr_reg[2]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(352[27:47])
    defparam round_ctr_reg_912__i2.GSR = "ENABLED";
    FD1P3IX round_ctr_reg_912__i1 (.D(n3[1]), .SP(round_ctr_we), .CD(n6361[2]), 
            .CK(clk_c), .Q(round_ctr_reg[1]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(352[27:47])
    defparam round_ctr_reg_912__i1.GSR = "ENABLED";
    LUT4 mux_17_i123_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [122]), 
         .D(key_mem_new[122]), .Z(key_mem_0__127__N_5728[122])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i123_3_lut_4_lut.init = 16'hf1e0;
    FD1P3IX rcon_reg_i0_i6 (.D(\rcon_logic.tmp_rcon [6]), .SP(rcon_we), 
            .CD(n15086), .CK(clk_c), .Q(\rcon_logic.tmp_rcon [7])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam rcon_reg_i0_i6.GSR = "ENABLED";
    FD1P3IX rcon_reg_i0_i5 (.D(\rcon_logic.tmp_rcon [5]), .SP(rcon_we), 
            .CD(n15086), .CK(clk_c), .Q(\rcon_logic.tmp_rcon [6])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam rcon_reg_i0_i5.GSR = "ENABLED";
    FD1P3IX rcon_reg_i0_i4 (.D(\rcon_logic.tmp_rcon [4]), .SP(rcon_we), 
            .CD(n15086), .CK(clk_c), .Q(\rcon_logic.tmp_rcon [5])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam rcon_reg_i0_i4.GSR = "ENABLED";
    FD1P3IX rcon_reg_i0_i1 (.D(\rcon_logic.tmp_rcon [1]), .SP(rcon_we), 
            .CD(n15086), .CK(clk_c), .Q(\rcon_logic.tmp_rcon [2])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(146[9] 167[12])
    defparam rcon_reg_i0_i1.GSR = "ENABLED";
    LUT4 mux_17_i124_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [123]), 
         .D(key_mem_new[123]), .Z(key_mem_0__127__N_5728[123])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i124_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i125_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [124]), 
         .D(key_mem_new[124]), .Z(key_mem_0__127__N_5728[124])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i125_3_lut_4_lut.init = 16'hf1e0;
    FD1P3IX round_ctr_reg_912__i0 (.D(n1_adj_9290), .SP(round_ctr_we), .CD(n6361[2]), 
            .CK(clk_c), .Q(round_ctr_reg[0]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(352[27:47])
    defparam round_ctr_reg_912__i0.GSR = "ENABLED";
    LUT4 mux_17_i126_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [125]), 
         .D(key_mem_new[125]), .Z(key_mem_0__127__N_5728[125])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i126_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i127_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [126]), 
         .D(key_mem_new[126]), .Z(key_mem_0__127__N_5728[126])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i127_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_17_i128_3_lut_4_lut (.A(n33912), .B(n33916), .C(\key_mem[6] [127]), 
         .D(key_mem_new[127]), .Z(key_mem_0__127__N_5728[127])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_17_i128_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_16_i1_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [0]), 
         .D(key_mem_new[0]), .Z(key_mem_0__127__N_5856[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i1_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i2_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [1]), 
         .D(key_mem_new[1]), .Z(key_mem_0__127__N_5856[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i2_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i3_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [2]), 
         .D(key_mem_new[2]), .Z(key_mem_0__127__N_5856[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i3_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25058 (.BLUT(n1_adj_9136), .ALUT(n2_adj_9135), .C0(\muxed_round_nr[1] ), 
          .Z(n30217));
    LUT4 mux_16_i4_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [3]), 
         .D(key_mem_new[3]), .Z(key_mem_0__127__N_5856[3])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i4_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i5_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [4]), 
         .D(key_mem_new[4]), .Z(key_mem_0__127__N_5856[4])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i5_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i6_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [5]), 
         .D(key_mem_new[5]), .Z(key_mem_0__127__N_5856[5])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i6_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25059 (.BLUT(n4_adj_9134), .ALUT(n5_adj_9133), .C0(\muxed_round_nr[1] ), 
          .Z(n30218));
    PFUMX i25060 (.BLUT(n8_adj_9132), .ALUT(n9_adj_9131), .C0(\muxed_round_nr[1] ), 
          .Z(n30219));
    LUT4 mux_16_i7_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [6]), 
         .D(key_mem_new[6]), .Z(key_mem_0__127__N_5856[6])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i7_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i8_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [7]), 
         .D(key_mem_new[7]), .Z(key_mem_0__127__N_5856[7])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i8_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i9_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [8]), 
         .D(key_mem_new[8]), .Z(key_mem_0__127__N_5856[8])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i9_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i10_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [9]), 
         .D(key_mem_new[9]), .Z(key_mem_0__127__N_5856[9])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i10_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i11_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [10]), 
         .D(key_mem_new[10]), .Z(key_mem_0__127__N_5856[10])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i11_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i12_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [11]), 
         .D(key_mem_new[11]), .Z(key_mem_0__127__N_5856[11])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i12_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i13_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [12]), 
         .D(key_mem_new[12]), .Z(key_mem_0__127__N_5856[12])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i13_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i14_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [13]), 
         .D(key_mem_new[13]), .Z(key_mem_0__127__N_5856[13])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i14_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i15_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [14]), 
         .D(key_mem_new[14]), .Z(key_mem_0__127__N_5856[14])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i15_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i16_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [15]), 
         .D(key_mem_new[15]), .Z(key_mem_0__127__N_5856[15])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i16_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i17_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [16]), 
         .D(key_mem_new[16]), .Z(key_mem_0__127__N_5856[16])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i17_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i18_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [17]), 
         .D(key_mem_new[17]), .Z(key_mem_0__127__N_5856[17])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i18_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i19_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [18]), 
         .D(key_mem_new[18]), .Z(key_mem_0__127__N_5856[18])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i19_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i20_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [19]), 
         .D(key_mem_new[19]), .Z(key_mem_0__127__N_5856[19])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i20_3_lut_4_lut.init = 16'hf2d0;
    FD1P3IX round_ctr_reg_912__i0_rep_649 (.D(n1_adj_9290), .SP(round_ctr_we), 
            .CD(n6361[2]), .CK(clk_c), .Q(n35834));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(352[27:47])
    defparam round_ctr_reg_912__i0_rep_649.GSR = "ENABLED";
    LUT4 mux_16_i21_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [20]), 
         .D(key_mem_new[20]), .Z(key_mem_0__127__N_5856[20])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i21_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i22_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [21]), 
         .D(key_mem_new[21]), .Z(key_mem_0__127__N_5856[21])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i22_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25725 (.BLUT(n8_adj_9127), .ALUT(n9_adj_9124), .C0(\muxed_round_nr[1] ), 
          .Z(n30884));
    PFUMX i25065 (.BLUT(n1_adj_9128), .ALUT(n2_adj_9126), .C0(\muxed_round_nr[1] ), 
          .Z(n30224));
    LUT4 mux_16_i23_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [22]), 
         .D(key_mem_new[22]), .Z(key_mem_0__127__N_5856[22])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i23_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i24_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [23]), 
         .D(key_mem_new[23]), .Z(key_mem_0__127__N_5856[23])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i24_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i25_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [24]), 
         .D(key_mem_new[24]), .Z(key_mem_0__127__N_5856[24])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i25_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i26_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [25]), 
         .D(key_mem_new[25]), .Z(key_mem_0__127__N_5856[25])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i26_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i27_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [26]), 
         .D(key_mem_new[26]), .Z(key_mem_0__127__N_5856[26])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i27_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i28_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [27]), 
         .D(key_mem_new[27]), .Z(key_mem_0__127__N_5856[27])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i28_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i29_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [28]), 
         .D(key_mem_new[28]), .Z(key_mem_0__127__N_5856[28])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i29_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i30_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [29]), 
         .D(key_mem_new[29]), .Z(key_mem_0__127__N_5856[29])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i30_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i31_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [30]), 
         .D(key_mem_new[30]), .Z(key_mem_0__127__N_5856[30])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i31_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i32_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [31]), 
         .D(key_mem_new[31]), .Z(key_mem_0__127__N_5856[31])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i32_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25066 (.BLUT(n4_adj_9125), .ALUT(n5_adj_9123), .C0(\muxed_round_nr[1] ), 
          .Z(n30225));
    LUT4 mux_16_i33_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [32]), 
         .D(key_mem_new[32]), .Z(key_mem_0__127__N_5856[32])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i33_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i34_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [33]), 
         .D(key_mem_new[33]), .Z(key_mem_0__127__N_5856[33])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i34_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25067 (.BLUT(n8_adj_9121), .ALUT(n9_adj_9118), .C0(\muxed_round_nr[1] ), 
          .Z(n30226));
    LUT4 mux_16_i35_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [34]), 
         .D(key_mem_new[34]), .Z(key_mem_0__127__N_5856[34])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i35_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i36_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [35]), 
         .D(key_mem_new[35]), .Z(key_mem_0__127__N_5856[35])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i36_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i37_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [36]), 
         .D(key_mem_new[36]), .Z(key_mem_0__127__N_5856[36])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i37_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i38_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [37]), 
         .D(key_mem_new[37]), .Z(key_mem_0__127__N_5856[37])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i38_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i39_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [38]), 
         .D(key_mem_new[38]), .Z(key_mem_0__127__N_5856[38])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i39_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i40_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [39]), 
         .D(key_mem_new[39]), .Z(key_mem_0__127__N_5856[39])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i40_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i41_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [40]), 
         .D(key_mem_new[40]), .Z(key_mem_0__127__N_5856[40])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i41_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i42_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [41]), 
         .D(key_mem_new[41]), .Z(key_mem_0__127__N_5856[41])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i42_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i43_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [42]), 
         .D(key_mem_new[42]), .Z(key_mem_0__127__N_5856[42])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i43_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i44_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [43]), 
         .D(key_mem_new[43]), .Z(key_mem_0__127__N_5856[43])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i44_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i45_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [44]), 
         .D(key_mem_new[44]), .Z(key_mem_0__127__N_5856[44])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i45_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i46_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [45]), 
         .D(key_mem_new[45]), .Z(key_mem_0__127__N_5856[45])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i46_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i47_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [46]), 
         .D(key_mem_new[46]), .Z(key_mem_0__127__N_5856[46])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i47_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i48_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [47]), 
         .D(key_mem_new[47]), .Z(key_mem_0__127__N_5856[47])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i48_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i49_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [48]), 
         .D(key_mem_new[48]), .Z(key_mem_0__127__N_5856[48])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i49_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i50_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [49]), 
         .D(key_mem_new[49]), .Z(key_mem_0__127__N_5856[49])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i50_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i51_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [50]), 
         .D(key_mem_new[50]), .Z(key_mem_0__127__N_5856[50])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i51_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i52_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [51]), 
         .D(key_mem_new[51]), .Z(key_mem_0__127__N_5856[51])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i52_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i53_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [52]), 
         .D(key_mem_new[52]), .Z(key_mem_0__127__N_5856[52])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i53_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i54_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [53]), 
         .D(key_mem_new[53]), .Z(key_mem_0__127__N_5856[53])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i54_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i55_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [54]), 
         .D(key_mem_new[54]), .Z(key_mem_0__127__N_5856[54])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i55_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i56_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [55]), 
         .D(key_mem_new[55]), .Z(key_mem_0__127__N_5856[55])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i56_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i57_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [56]), 
         .D(key_mem_new[56]), .Z(key_mem_0__127__N_5856[56])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i57_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i58_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [57]), 
         .D(key_mem_new[57]), .Z(key_mem_0__127__N_5856[57])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i58_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i59_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [58]), 
         .D(key_mem_new[58]), .Z(key_mem_0__127__N_5856[58])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i59_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i60_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [59]), 
         .D(key_mem_new[59]), .Z(key_mem_0__127__N_5856[59])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i60_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i61_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [60]), 
         .D(key_mem_new[60]), .Z(key_mem_0__127__N_5856[60])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i61_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i62_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [61]), 
         .D(key_mem_new[61]), .Z(key_mem_0__127__N_5856[61])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i62_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i63_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [62]), 
         .D(key_mem_new[62]), .Z(key_mem_0__127__N_5856[62])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i63_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i64_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [63]), 
         .D(key_mem_new[63]), .Z(key_mem_0__127__N_5856[63])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i64_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25730 (.BLUT(n1_adj_9120), .ALUT(n2_adj_9119), .C0(\muxed_round_nr[1] ), 
          .Z(n30889));
    LUT4 mux_16_i65_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [64]), 
         .D(key_mem_new[64]), .Z(key_mem_0__127__N_5856[64])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i65_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i66_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [65]), 
         .D(key_mem_new[65]), .Z(key_mem_0__127__N_5856[65])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i66_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i67_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [66]), 
         .D(key_mem_new[66]), .Z(key_mem_0__127__N_5856[66])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i67_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i68_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [67]), 
         .D(key_mem_new[67]), .Z(key_mem_0__127__N_5856[67])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i68_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i69_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [68]), 
         .D(key_mem_new[68]), .Z(key_mem_0__127__N_5856[68])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i69_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i70_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [69]), 
         .D(key_mem_new[69]), .Z(key_mem_0__127__N_5856[69])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i70_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i71_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [70]), 
         .D(key_mem_new[70]), .Z(key_mem_0__127__N_5856[70])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i71_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i72_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [71]), 
         .D(key_mem_new[71]), .Z(key_mem_0__127__N_5856[71])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i72_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25731 (.BLUT(n4_adj_9116), .ALUT(n5_adj_9115), .C0(\muxed_round_nr[1] ), 
          .Z(n30890));
    LUT4 mux_16_i73_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [72]), 
         .D(key_mem_new[72]), .Z(key_mem_0__127__N_5856[72])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i73_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i74_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [73]), 
         .D(key_mem_new[73]), .Z(key_mem_0__127__N_5856[73])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i74_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i75_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [74]), 
         .D(key_mem_new[74]), .Z(key_mem_0__127__N_5856[74])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i75_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i76_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [75]), 
         .D(key_mem_new[75]), .Z(key_mem_0__127__N_5856[75])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i76_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25072 (.BLUT(n1_adj_9114), .ALUT(n2_adj_9113), .C0(\muxed_round_nr[1] ), 
          .Z(n30231));
    LUT4 mux_16_i77_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [76]), 
         .D(key_mem_new[76]), .Z(key_mem_0__127__N_5856[76])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i77_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i78_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [77]), 
         .D(key_mem_new[77]), .Z(key_mem_0__127__N_5856[77])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i78_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i79_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [78]), 
         .D(key_mem_new[78]), .Z(key_mem_0__127__N_5856[78])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i79_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i80_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [79]), 
         .D(key_mem_new[79]), .Z(key_mem_0__127__N_5856[79])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i80_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i81_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [80]), 
         .D(key_mem_new[80]), .Z(key_mem_0__127__N_5856[80])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i81_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25073 (.BLUT(n4_adj_9112), .ALUT(n5_adj_9111), .C0(\muxed_round_nr[1] ), 
          .Z(n30232));
    LUT4 mux_16_i82_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [81]), 
         .D(key_mem_new[81]), .Z(key_mem_0__127__N_5856[81])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i82_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i83_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [82]), 
         .D(key_mem_new[82]), .Z(key_mem_0__127__N_5856[82])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i83_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25074 (.BLUT(n8_adj_9110), .ALUT(n9_adj_9109), .C0(\muxed_round_nr[1] ), 
          .Z(n30233));
    LUT4 mux_16_i84_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [83]), 
         .D(key_mem_new[83]), .Z(key_mem_0__127__N_5856[83])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i84_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i85_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [84]), 
         .D(key_mem_new[84]), .Z(key_mem_0__127__N_5856[84])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i85_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i86_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [85]), 
         .D(key_mem_new[85]), .Z(key_mem_0__127__N_5856[85])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i86_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i87_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [86]), 
         .D(key_mem_new[86]), .Z(key_mem_0__127__N_5856[86])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i87_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i88_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [87]), 
         .D(key_mem_new[87]), .Z(key_mem_0__127__N_5856[87])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i88_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i89_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [88]), 
         .D(key_mem_new[88]), .Z(key_mem_0__127__N_5856[88])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i89_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i90_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [89]), 
         .D(key_mem_new[89]), .Z(key_mem_0__127__N_5856[89])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i90_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i91_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [90]), 
         .D(key_mem_new[90]), .Z(key_mem_0__127__N_5856[90])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i91_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i92_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [91]), 
         .D(key_mem_new[91]), .Z(key_mem_0__127__N_5856[91])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i92_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i93_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [92]), 
         .D(key_mem_new[92]), .Z(key_mem_0__127__N_5856[92])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i93_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i94_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [93]), 
         .D(key_mem_new[93]), .Z(key_mem_0__127__N_5856[93])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i94_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i95_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [94]), 
         .D(key_mem_new[94]), .Z(key_mem_0__127__N_5856[94])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i95_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i96_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [95]), 
         .D(key_mem_new[95]), .Z(key_mem_0__127__N_5856[95])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i96_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i97_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [96]), 
         .D(key_mem_new[96]), .Z(key_mem_0__127__N_5856[96])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i97_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i98_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [97]), 
         .D(key_mem_new[97]), .Z(key_mem_0__127__N_5856[97])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i98_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i99_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [98]), 
         .D(key_mem_new[98]), .Z(key_mem_0__127__N_5856[98])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i99_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i100_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [99]), 
         .D(key_mem_new[99]), .Z(key_mem_0__127__N_5856[99])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i100_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i101_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [100]), 
         .D(key_mem_new[100]), .Z(key_mem_0__127__N_5856[100])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i101_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i102_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [101]), 
         .D(key_mem_new[101]), .Z(key_mem_0__127__N_5856[101])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i102_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i103_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [102]), 
         .D(key_mem_new[102]), .Z(key_mem_0__127__N_5856[102])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i103_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i104_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [103]), 
         .D(key_mem_new[103]), .Z(key_mem_0__127__N_5856[103])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i104_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25079 (.BLUT(n1_adj_9107), .ALUT(n2_adj_9106), .C0(\muxed_round_nr[1] ), 
          .Z(n30238));
    LUT4 mux_16_i105_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [104]), 
         .D(key_mem_new[104]), .Z(key_mem_0__127__N_5856[104])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i105_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i106_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [105]), 
         .D(key_mem_new[105]), .Z(key_mem_0__127__N_5856[105])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i106_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i107_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [106]), 
         .D(key_mem_new[106]), .Z(key_mem_0__127__N_5856[106])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i107_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i108_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [107]), 
         .D(key_mem_new[107]), .Z(key_mem_0__127__N_5856[107])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i108_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i109_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [108]), 
         .D(key_mem_new[108]), .Z(key_mem_0__127__N_5856[108])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i109_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i110_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [109]), 
         .D(key_mem_new[109]), .Z(key_mem_0__127__N_5856[109])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i110_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i111_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [110]), 
         .D(key_mem_new[110]), .Z(key_mem_0__127__N_5856[110])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i111_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i112_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [111]), 
         .D(key_mem_new[111]), .Z(key_mem_0__127__N_5856[111])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i112_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i113_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [112]), 
         .D(key_mem_new[112]), .Z(key_mem_0__127__N_5856[112])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i113_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25080 (.BLUT(n4_adj_9105), .ALUT(n5_adj_9104), .C0(\muxed_round_nr[1] ), 
          .Z(n30239));
    LUT4 mux_16_i114_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [113]), 
         .D(key_mem_new[113]), .Z(key_mem_0__127__N_5856[113])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i114_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25732 (.BLUT(n8_adj_9093), .ALUT(n9_adj_9092), .C0(\muxed_round_nr[1] ), 
          .Z(n30891));
    LUT4 mux_16_i115_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [114]), 
         .D(key_mem_new[114]), .Z(key_mem_0__127__N_5856[114])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i115_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i116_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [115]), 
         .D(key_mem_new[115]), .Z(key_mem_0__127__N_5856[115])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i116_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i117_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [116]), 
         .D(key_mem_new[116]), .Z(key_mem_0__127__N_5856[116])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i117_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i118_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [117]), 
         .D(key_mem_new[117]), .Z(key_mem_0__127__N_5856[117])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i118_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i119_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [118]), 
         .D(key_mem_new[118]), .Z(key_mem_0__127__N_5856[118])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i119_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i120_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [119]), 
         .D(key_mem_new[119]), .Z(key_mem_0__127__N_5856[119])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i120_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i121_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [120]), 
         .D(key_mem_new[120]), .Z(key_mem_0__127__N_5856[120])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i121_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i122_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [121]), 
         .D(key_mem_new[121]), .Z(key_mem_0__127__N_5856[121])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i122_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25081 (.BLUT(n8_adj_9103), .ALUT(n9_adj_9102), .C0(\muxed_round_nr[1] ), 
          .Z(n30240));
    LUT4 mux_16_i123_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [122]), 
         .D(key_mem_new[122]), .Z(key_mem_0__127__N_5856[122])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i123_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i124_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [123]), 
         .D(key_mem_new[123]), .Z(key_mem_0__127__N_5856[123])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i124_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i125_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [124]), 
         .D(key_mem_new[124]), .Z(key_mem_0__127__N_5856[124])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i125_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i126_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [125]), 
         .D(key_mem_new[125]), .Z(key_mem_0__127__N_5856[125])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i126_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i127_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [126]), 
         .D(key_mem_new[126]), .Z(key_mem_0__127__N_5856[126])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i127_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_16_i128_3_lut_4_lut (.A(n33938), .B(n33916), .C(\key_mem[7] [127]), 
         .D(key_mem_new[127]), .Z(key_mem_0__127__N_5856[127])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_16_i128_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_15_i65_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [64]), 
         .D(key_mem_new[64]), .Z(key_mem_0__127__N_5984[64])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i65_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i39_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [38]), 
         .D(key_mem_new[38]), .Z(key_mem_0__127__N_5984[38])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i39_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i40_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [39]), 
         .D(key_mem_new[39]), .Z(key_mem_0__127__N_5984[39])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i40_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i41_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [40]), 
         .D(key_mem_new[40]), .Z(key_mem_0__127__N_5984[40])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i41_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i42_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [41]), 
         .D(key_mem_new[41]), .Z(key_mem_0__127__N_5984[41])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i42_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i43_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [42]), 
         .D(key_mem_new[42]), .Z(key_mem_0__127__N_5984[42])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i43_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i44_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [43]), 
         .D(key_mem_new[43]), .Z(key_mem_0__127__N_5984[43])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i44_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i45_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [44]), 
         .D(key_mem_new[44]), .Z(key_mem_0__127__N_5984[44])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i45_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i46_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [45]), 
         .D(key_mem_new[45]), .Z(key_mem_0__127__N_5984[45])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i46_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i47_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [46]), 
         .D(key_mem_new[46]), .Z(key_mem_0__127__N_5984[46])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i47_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i48_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [47]), 
         .D(key_mem_new[47]), .Z(key_mem_0__127__N_5984[47])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i48_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i49_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [48]), 
         .D(key_mem_new[48]), .Z(key_mem_0__127__N_5984[48])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i49_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i50_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [49]), 
         .D(key_mem_new[49]), .Z(key_mem_0__127__N_5984[49])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i50_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i51_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [50]), 
         .D(key_mem_new[50]), .Z(key_mem_0__127__N_5984[50])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i51_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i52_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [51]), 
         .D(key_mem_new[51]), .Z(key_mem_0__127__N_5984[51])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i52_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25086 (.BLUT(n1_adj_9100), .ALUT(n2_adj_9099), .C0(\muxed_round_nr[1] ), 
          .Z(n30245));
    LUT4 mux_15_i53_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [52]), 
         .D(key_mem_new[52]), .Z(key_mem_0__127__N_5984[52])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i53_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i54_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [53]), 
         .D(key_mem_new[53]), .Z(key_mem_0__127__N_5984[53])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i54_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25087 (.BLUT(n4_adj_9098), .ALUT(n5_adj_9097), .C0(\muxed_round_nr[1] ), 
          .Z(n30246));
    LUT4 mux_15_i55_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [54]), 
         .D(key_mem_new[54]), .Z(key_mem_0__127__N_5984[54])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i55_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i56_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [55]), 
         .D(key_mem_new[55]), .Z(key_mem_0__127__N_5984[55])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i56_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i57_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [56]), 
         .D(key_mem_new[56]), .Z(key_mem_0__127__N_5984[56])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i57_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25088 (.BLUT(n8_adj_9096), .ALUT(n9_adj_9095), .C0(\muxed_round_nr[1] ), 
          .Z(n30247));
    LUT4 mux_15_i58_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [57]), 
         .D(key_mem_new[57]), .Z(key_mem_0__127__N_5984[57])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i58_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i59_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [58]), 
         .D(key_mem_new[58]), .Z(key_mem_0__127__N_5984[58])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i59_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i60_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [59]), 
         .D(key_mem_new[59]), .Z(key_mem_0__127__N_5984[59])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i60_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i61_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [60]), 
         .D(key_mem_new[60]), .Z(key_mem_0__127__N_5984[60])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i61_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i62_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [61]), 
         .D(key_mem_new[61]), .Z(key_mem_0__127__N_5984[61])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i62_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i63_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [62]), 
         .D(key_mem_new[62]), .Z(key_mem_0__127__N_5984[62])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i63_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i64_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [63]), 
         .D(key_mem_new[63]), .Z(key_mem_0__127__N_5984[63])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i64_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i1_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [0]), 
         .D(key_mem_new[0]), .Z(key_mem_0__127__N_5984[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i2_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [1]), 
         .D(key_mem_new[1]), .Z(key_mem_0__127__N_5984[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i3_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [2]), 
         .D(key_mem_new[2]), .Z(key_mem_0__127__N_5984[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i4_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [3]), 
         .D(key_mem_new[3]), .Z(key_mem_0__127__N_5984[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i5_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [4]), 
         .D(key_mem_new[4]), .Z(key_mem_0__127__N_5984[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i6_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [5]), 
         .D(key_mem_new[5]), .Z(key_mem_0__127__N_5984[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i7_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [6]), 
         .D(key_mem_new[6]), .Z(key_mem_0__127__N_5984[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i8_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [7]), 
         .D(key_mem_new[7]), .Z(key_mem_0__127__N_5984[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i9_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [8]), 
         .D(key_mem_new[8]), .Z(key_mem_0__127__N_5984[8])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i9_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i10_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [9]), 
         .D(key_mem_new[9]), .Z(key_mem_0__127__N_5984[9])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i10_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i11_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [10]), 
         .D(key_mem_new[10]), .Z(key_mem_0__127__N_5984[10])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i11_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i12_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [11]), 
         .D(key_mem_new[11]), .Z(key_mem_0__127__N_5984[11])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i12_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i13_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [12]), 
         .D(key_mem_new[12]), .Z(key_mem_0__127__N_5984[12])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i13_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i14_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [13]), 
         .D(key_mem_new[13]), .Z(key_mem_0__127__N_5984[13])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i14_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25093 (.BLUT(n1_adj_9091), .ALUT(n2_adj_9089), .C0(\muxed_round_nr[1] ), 
          .Z(n30252));
    LUT4 mux_15_i15_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [14]), 
         .D(key_mem_new[14]), .Z(key_mem_0__127__N_5984[14])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i15_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i16_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [15]), 
         .D(key_mem_new[15]), .Z(key_mem_0__127__N_5984[15])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i16_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i17_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [16]), 
         .D(key_mem_new[16]), .Z(key_mem_0__127__N_5984[16])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i17_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i18_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [17]), 
         .D(key_mem_new[17]), .Z(key_mem_0__127__N_5984[17])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i18_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i19_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [18]), 
         .D(key_mem_new[18]), .Z(key_mem_0__127__N_5984[18])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i19_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i20_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [19]), 
         .D(key_mem_new[19]), .Z(key_mem_0__127__N_5984[19])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i20_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i21_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [20]), 
         .D(key_mem_new[20]), .Z(key_mem_0__127__N_5984[20])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i21_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i22_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [21]), 
         .D(key_mem_new[21]), .Z(key_mem_0__127__N_5984[21])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i22_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i23_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [22]), 
         .D(key_mem_new[22]), .Z(key_mem_0__127__N_5984[22])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i23_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i24_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [23]), 
         .D(key_mem_new[23]), .Z(key_mem_0__127__N_5984[23])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i24_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i25_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [24]), 
         .D(key_mem_new[24]), .Z(key_mem_0__127__N_5984[24])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i25_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i26_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [25]), 
         .D(key_mem_new[25]), .Z(key_mem_0__127__N_5984[25])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i26_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i27_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [26]), 
         .D(key_mem_new[26]), .Z(key_mem_0__127__N_5984[26])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i27_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i28_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [27]), 
         .D(key_mem_new[27]), .Z(key_mem_0__127__N_5984[27])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i28_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i29_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [28]), 
         .D(key_mem_new[28]), .Z(key_mem_0__127__N_5984[28])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i29_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i30_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [29]), 
         .D(key_mem_new[29]), .Z(key_mem_0__127__N_5984[29])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i30_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i31_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [30]), 
         .D(key_mem_new[30]), .Z(key_mem_0__127__N_5984[30])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i31_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i32_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [31]), 
         .D(key_mem_new[31]), .Z(key_mem_0__127__N_5984[31])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i32_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i33_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [32]), 
         .D(key_mem_new[32]), .Z(key_mem_0__127__N_5984[32])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i33_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i34_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [33]), 
         .D(key_mem_new[33]), .Z(key_mem_0__127__N_5984[33])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i34_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i35_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [34]), 
         .D(key_mem_new[34]), .Z(key_mem_0__127__N_5984[34])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i35_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i36_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [35]), 
         .D(key_mem_new[35]), .Z(key_mem_0__127__N_5984[35])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i36_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i37_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [36]), 
         .D(key_mem_new[36]), .Z(key_mem_0__127__N_5984[36])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i37_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i38_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [37]), 
         .D(key_mem_new[37]), .Z(key_mem_0__127__N_5984[37])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i38_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i66_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [65]), 
         .D(key_mem_new[65]), .Z(key_mem_0__127__N_5984[65])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i66_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i67_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [66]), 
         .D(key_mem_new[66]), .Z(key_mem_0__127__N_5984[66])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i67_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i68_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [67]), 
         .D(key_mem_new[67]), .Z(key_mem_0__127__N_5984[67])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i68_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i69_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [68]), 
         .D(key_mem_new[68]), .Z(key_mem_0__127__N_5984[68])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i69_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i70_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [69]), 
         .D(key_mem_new[69]), .Z(key_mem_0__127__N_5984[69])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i70_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i71_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [70]), 
         .D(key_mem_new[70]), .Z(key_mem_0__127__N_5984[70])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i71_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i72_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [71]), 
         .D(key_mem_new[71]), .Z(key_mem_0__127__N_5984[71])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i72_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i73_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [72]), 
         .D(key_mem_new[72]), .Z(key_mem_0__127__N_5984[72])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i73_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i74_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [73]), 
         .D(key_mem_new[73]), .Z(key_mem_0__127__N_5984[73])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i74_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i75_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [74]), 
         .D(key_mem_new[74]), .Z(key_mem_0__127__N_5984[74])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i75_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i76_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [75]), 
         .D(key_mem_new[75]), .Z(key_mem_0__127__N_5984[75])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i76_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i77_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [76]), 
         .D(key_mem_new[76]), .Z(key_mem_0__127__N_5984[76])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i77_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i78_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [77]), 
         .D(key_mem_new[77]), .Z(key_mem_0__127__N_5984[77])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i78_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i79_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [78]), 
         .D(key_mem_new[78]), .Z(key_mem_0__127__N_5984[78])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i79_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i80_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [79]), 
         .D(key_mem_new[79]), .Z(key_mem_0__127__N_5984[79])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i80_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i81_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [80]), 
         .D(key_mem_new[80]), .Z(key_mem_0__127__N_5984[80])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i81_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i82_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [81]), 
         .D(key_mem_new[81]), .Z(key_mem_0__127__N_5984[81])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i82_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i83_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [82]), 
         .D(key_mem_new[82]), .Z(key_mem_0__127__N_5984[82])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i83_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i84_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [83]), 
         .D(key_mem_new[83]), .Z(key_mem_0__127__N_5984[83])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i84_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i85_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [84]), 
         .D(key_mem_new[84]), .Z(key_mem_0__127__N_5984[84])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i85_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i86_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [85]), 
         .D(key_mem_new[85]), .Z(key_mem_0__127__N_5984[85])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i86_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i87_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [86]), 
         .D(key_mem_new[86]), .Z(key_mem_0__127__N_5984[86])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i87_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i88_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [87]), 
         .D(key_mem_new[87]), .Z(key_mem_0__127__N_5984[87])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i88_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i89_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [88]), 
         .D(key_mem_new[88]), .Z(key_mem_0__127__N_5984[88])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i89_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i90_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [89]), 
         .D(key_mem_new[89]), .Z(key_mem_0__127__N_5984[89])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i90_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i91_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [90]), 
         .D(key_mem_new[90]), .Z(key_mem_0__127__N_5984[90])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i91_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i92_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [91]), 
         .D(key_mem_new[91]), .Z(key_mem_0__127__N_5984[91])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i92_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25094 (.BLUT(n4_adj_9088), .ALUT(n5_adj_9087), .C0(\muxed_round_nr[1] ), 
          .Z(n30253));
    LUT4 mux_15_i93_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [92]), 
         .D(key_mem_new[92]), .Z(key_mem_0__127__N_5984[92])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i93_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i94_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [93]), 
         .D(key_mem_new[93]), .Z(key_mem_0__127__N_5984[93])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i94_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i95_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [94]), 
         .D(key_mem_new[94]), .Z(key_mem_0__127__N_5984[94])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i95_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i96_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [95]), 
         .D(key_mem_new[95]), .Z(key_mem_0__127__N_5984[95])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i96_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25095 (.BLUT(n8_adj_9086), .ALUT(n9_adj_9085), .C0(\muxed_round_nr[1] ), 
          .Z(n30254));
    LUT4 mux_15_i97_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [96]), 
         .D(key_mem_new[96]), .Z(key_mem_0__127__N_5984[96])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i97_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i11220 (.BLUT(n16797), .ALUT(n16802), .C0(n35835), .Z(n16803));
    LUT4 mux_15_i98_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [97]), 
         .D(key_mem_new[97]), .Z(key_mem_0__127__N_5984[97])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i98_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i99_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [98]), 
         .D(key_mem_new[98]), .Z(key_mem_0__127__N_5984[98])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i99_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i100_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [99]), 
         .D(key_mem_new[99]), .Z(key_mem_0__127__N_5984[99])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i100_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i101_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [100]), 
         .D(key_mem_new[100]), .Z(key_mem_0__127__N_5984[100])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i101_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i102_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [101]), 
         .D(key_mem_new[101]), .Z(key_mem_0__127__N_5984[101])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i102_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i103_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [102]), 
         .D(key_mem_new[102]), .Z(key_mem_0__127__N_5984[102])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i103_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i104_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [103]), 
         .D(key_mem_new[103]), .Z(key_mem_0__127__N_5984[103])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i104_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i105_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [104]), 
         .D(key_mem_new[104]), .Z(key_mem_0__127__N_5984[104])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i105_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i106_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [105]), 
         .D(key_mem_new[105]), .Z(key_mem_0__127__N_5984[105])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i106_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i107_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [106]), 
         .D(key_mem_new[106]), .Z(key_mem_0__127__N_5984[106])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i107_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i108_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [107]), 
         .D(key_mem_new[107]), .Z(key_mem_0__127__N_5984[107])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i108_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i109_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [108]), 
         .D(key_mem_new[108]), .Z(key_mem_0__127__N_5984[108])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i109_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i110_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [109]), 
         .D(key_mem_new[109]), .Z(key_mem_0__127__N_5984[109])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i110_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i111_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [110]), 
         .D(key_mem_new[110]), .Z(key_mem_0__127__N_5984[110])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i111_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i112_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [111]), 
         .D(key_mem_new[111]), .Z(key_mem_0__127__N_5984[111])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i112_3_lut_4_lut.init = 16'hf1e0;
    PFUMX keylen_I_0_Mux_95_i1 (.BLUT(key_mem_new_127__N_7264[95]), .ALUT(prev_key1_new_127__N_7520[95]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[95])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    LUT4 mux_15_i113_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [112]), 
         .D(key_mem_new[112]), .Z(key_mem_0__127__N_5984[112])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i113_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i114_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [113]), 
         .D(key_mem_new[113]), .Z(key_mem_0__127__N_5984[113])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i114_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25100 (.BLUT(n1_adj_9082), .ALUT(n2_adj_9081), .C0(\muxed_round_nr[1] ), 
          .Z(n30259));
    LUT4 mux_15_i115_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [114]), 
         .D(key_mem_new[114]), .Z(key_mem_0__127__N_5984[114])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i115_3_lut_4_lut.init = 16'hf1e0;
    PFUMX keylen_I_0_Mux_94_i1 (.BLUT(key_mem_new_127__N_7264[94]), .ALUT(prev_key1_new_127__N_7520[94]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[94])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    LUT4 mux_15_i116_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [115]), 
         .D(key_mem_new[115]), .Z(key_mem_0__127__N_5984[115])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i116_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i117_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [116]), 
         .D(key_mem_new[116]), .Z(key_mem_0__127__N_5984[116])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i117_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i118_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [117]), 
         .D(key_mem_new[117]), .Z(key_mem_0__127__N_5984[117])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i118_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25737 (.BLUT(n1_adj_9080), .ALUT(n2_adj_9078), .C0(\muxed_round_nr[1] ), 
          .Z(n30896));
    FD1P3AX key_mem_ctrl_reg_FSM_i0_i1 (.D(n6361[2]), .SP(key_mem_ctrl_we), 
            .CK(clk_c), .Q(n6361[1]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam key_mem_ctrl_reg_FSM_i0_i1.GSR = "ENABLED";
    LUT4 mux_15_i119_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [118]), 
         .D(key_mem_new[118]), .Z(key_mem_0__127__N_5984[118])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i119_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i120_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [119]), 
         .D(key_mem_new[119]), .Z(key_mem_0__127__N_5984[119])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i120_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i121_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [120]), 
         .D(key_mem_new[120]), .Z(key_mem_0__127__N_5984[120])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i121_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i122_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [121]), 
         .D(key_mem_new[121]), .Z(key_mem_0__127__N_5984[121])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i122_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i123_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [122]), 
         .D(key_mem_new[122]), .Z(key_mem_0__127__N_5984[122])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i123_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i124_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [123]), 
         .D(key_mem_new[123]), .Z(key_mem_0__127__N_5984[123])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i124_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i125_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [124]), 
         .D(key_mem_new[124]), .Z(key_mem_0__127__N_5984[124])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i125_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i126_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [125]), 
         .D(key_mem_new[125]), .Z(key_mem_0__127__N_5984[125])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i126_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i127_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [126]), 
         .D(key_mem_new[126]), .Z(key_mem_0__127__N_5984[126])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i127_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_15_i128_3_lut_4_lut (.A(n33943), .B(n33937), .C(\key_mem[8] [127]), 
         .D(key_mem_new[127]), .Z(key_mem_0__127__N_5984[127])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_15_i128_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25101 (.BLUT(n4_adj_9079), .ALUT(n5_adj_9077), .C0(\muxed_round_nr[1] ), 
          .Z(n30260));
    PFUMX keylen_I_0_Mux_93_i1 (.BLUT(key_mem_new_127__N_7264[93]), .ALUT(prev_key1_new_127__N_7520[93]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[93])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    PFUMX i25102 (.BLUT(n8_adj_9076), .ALUT(n9_adj_9075), .C0(\muxed_round_nr[1] ), 
          .Z(n30261));
    PFUMX keylen_I_0_Mux_92_i1 (.BLUT(key_mem_new_127__N_7264[92]), .ALUT(prev_key1_new_127__N_7520[92]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[92])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    PFUMX keylen_I_0_Mux_91_i1 (.BLUT(key_mem_new_127__N_7264[91]), .ALUT(prev_key1_new_127__N_7520[91]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[91])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    PFUMX i25107 (.BLUT(n1_adj_9073), .ALUT(n2_adj_9072), .C0(\muxed_round_nr[1] ), 
          .Z(n30266));
    PFUMX keylen_I_0_Mux_90_i1 (.BLUT(key_mem_new_127__N_7264[90]), .ALUT(prev_key1_new_127__N_7520[90]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[90])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    PFUMX keylen_I_0_Mux_89_i1 (.BLUT(key_mem_new_127__N_7264[89]), .ALUT(prev_key1_new_127__N_7520[89]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[89])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    PFUMX i25108 (.BLUT(n4_adj_9071), .ALUT(n5_adj_9070), .C0(\muxed_round_nr[1] ), 
          .Z(n30267));
    PFUMX keylen_I_0_Mux_88_i1 (.BLUT(key_mem_new_127__N_7264[88]), .ALUT(prev_key1_new_127__N_7520[88]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[88])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    PFUMX i25109 (.BLUT(n8_adj_9069), .ALUT(n9_adj_9068), .C0(\muxed_round_nr[1] ), 
          .Z(n30268));
    PFUMX i11281 (.BLUT(n16857), .ALUT(n16862), .C0(n35835), .Z(n16863));
    PFUMX i11342 (.BLUT(n16917), .ALUT(n16922), .C0(n35835), .Z(n16923));
    PFUMX i25114 (.BLUT(n1_adj_9065), .ALUT(n2_adj_9063), .C0(\muxed_round_nr[1] ), 
          .Z(n30273));
    PFUMX i11403 (.BLUT(n16977), .ALUT(n16982), .C0(n35835), .Z(n16983));
    PFUMX i25115 (.BLUT(n4_adj_9062), .ALUT(n5_adj_9060), .C0(\muxed_round_nr[1] ), 
          .Z(n30274));
    PFUMX i25738 (.BLUT(n4_adj_9045), .ALUT(n5_adj_9044), .C0(\muxed_round_nr[1] ), 
          .Z(n30897));
    PFUMX i11464 (.BLUT(n17037), .ALUT(n17042), .C0(n35835), .Z(n17043));
    PFUMX i25116 (.BLUT(n8_adj_9058), .ALUT(n9_adj_9057), .C0(\muxed_round_nr[1] ), 
          .Z(n30275));
    PFUMX i11525 (.BLUT(n17097), .ALUT(n17102), .C0(n35835), .Z(n17103));
    PFUMX i11586 (.BLUT(n17157), .ALUT(n17162), .C0(n35835), .Z(n17163));
    PFUMX i25121 (.BLUT(n1_adj_9053), .ALUT(n2_adj_9052), .C0(\muxed_round_nr[1] ), 
          .Z(n30280));
    PFUMX i11647 (.BLUT(n17217), .ALUT(n17222), .C0(n35835), .Z(n17223));
    PFUMX i25122 (.BLUT(n4_adj_9050), .ALUT(n5_adj_9049), .C0(\muxed_round_nr[1] ), 
          .Z(n30281));
    PFUMX i9702 (.BLUT(n15304), .ALUT(n15309), .C0(n35835), .Z(n15310));
    PFUMX i25123 (.BLUT(n8_adj_9047), .ALUT(n9_adj_9043), .C0(\muxed_round_nr[1] ), 
          .Z(n30282));
    PFUMX i9817 (.BLUT(n15417), .ALUT(n15422), .C0(n35835), .Z(n15423));
    PFUMX i9878 (.BLUT(n15477), .ALUT(n15482), .C0(n35835), .Z(n15483));
    PFUMX i9939 (.BLUT(n15537), .ALUT(n15542), .C0(n35835), .Z(n15543));
    PFUMX i25128 (.BLUT(n1_adj_9039), .ALUT(n2_adj_9038), .C0(\muxed_round_nr[1] ), 
          .Z(n30287));
    PFUMX i25739 (.BLUT(n8_adj_9037), .ALUT(n9_adj_9036), .C0(\muxed_round_nr[1] ), 
          .Z(n30898));
    PFUMX i10000 (.BLUT(n15597), .ALUT(n15602), .C0(n35835), .Z(n15603));
    PFUMX i25129 (.BLUT(n4_adj_9035), .ALUT(n5_adj_9033), .C0(\muxed_round_nr[1] ), 
          .Z(n30288));
    PFUMX i10061 (.BLUT(n15657), .ALUT(n15662), .C0(n35835), .Z(n15663));
    LUT4 mux_14_i65_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [64]), 
         .D(key_mem_new[64]), .Z(key_mem_0__127__N_6112[64])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i65_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i39_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [38]), 
         .D(key_mem_new[38]), .Z(key_mem_0__127__N_6112[38])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i39_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i40_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [39]), 
         .D(key_mem_new[39]), .Z(key_mem_0__127__N_6112[39])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i40_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i38_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [37]), 
         .D(key_mem_new[37]), .Z(key_mem_0__127__N_6112[37])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i38_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25130 (.BLUT(n8_adj_9031), .ALUT(n9_adj_9030), .C0(\muxed_round_nr[1] ), 
          .Z(n30289));
    PFUMX i10122 (.BLUT(n15717), .ALUT(n15722), .C0(n35835), .Z(n15723));
    LUT4 mux_14_i42_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [41]), 
         .D(key_mem_new[41]), .Z(key_mem_0__127__N_6112[41])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i42_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i10183 (.BLUT(n15777), .ALUT(n15782), .C0(n35835), .Z(n15783));
    LUT4 mux_14_i41_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [40]), 
         .D(key_mem_new[40]), .Z(key_mem_0__127__N_6112[40])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i41_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25135 (.BLUT(n1_adj_9026), .ALUT(n2_adj_9025), .C0(\muxed_round_nr[1] ), 
          .Z(n30294));
    LUT4 mux_14_i44_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [43]), 
         .D(key_mem_new[43]), .Z(key_mem_0__127__N_6112[43])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i44_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i43_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [42]), 
         .D(key_mem_new[42]), .Z(key_mem_0__127__N_6112[42])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i43_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i46_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [45]), 
         .D(key_mem_new[45]), .Z(key_mem_0__127__N_6112[45])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i46_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i45_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [44]), 
         .D(key_mem_new[44]), .Z(key_mem_0__127__N_6112[44])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i45_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i48_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [47]), 
         .D(key_mem_new[47]), .Z(key_mem_0__127__N_6112[47])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i48_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i47_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [46]), 
         .D(key_mem_new[46]), .Z(key_mem_0__127__N_6112[46])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i47_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i10244 (.BLUT(n15837), .ALUT(n15842), .C0(n35835), .Z(n15843));
    LUT4 mux_14_i50_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [49]), 
         .D(key_mem_new[49]), .Z(key_mem_0__127__N_6112[49])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i50_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i49_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [48]), 
         .D(key_mem_new[48]), .Z(key_mem_0__127__N_6112[48])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i49_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i52_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [51]), 
         .D(key_mem_new[51]), .Z(key_mem_0__127__N_6112[51])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i52_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25136 (.BLUT(n4_adj_9023), .ALUT(n5_adj_9022), .C0(\muxed_round_nr[1] ), 
          .Z(n30295));
    PFUMX i10305 (.BLUT(n15897), .ALUT(n15902), .C0(n35835), .Z(n15903));
    LUT4 mux_14_i51_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [50]), 
         .D(key_mem_new[50]), .Z(key_mem_0__127__N_6112[50])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i51_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25137 (.BLUT(n8_adj_9018), .ALUT(n9_adj_9017), .C0(\muxed_round_nr[1] ), 
          .Z(n30296));
    LUT4 mux_14_i54_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [53]), 
         .D(key_mem_new[53]), .Z(key_mem_0__127__N_6112[53])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i54_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i10366 (.BLUT(n15957), .ALUT(n15962), .C0(n35835), .Z(n15963));
    LUT4 mux_14_i53_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [52]), 
         .D(key_mem_new[52]), .Z(key_mem_0__127__N_6112[52])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i53_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i56_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [55]), 
         .D(key_mem_new[55]), .Z(key_mem_0__127__N_6112[55])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i56_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i55_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [54]), 
         .D(key_mem_new[54]), .Z(key_mem_0__127__N_6112[54])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i55_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i58_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [57]), 
         .D(key_mem_new[57]), .Z(key_mem_0__127__N_6112[57])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i58_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i57_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [56]), 
         .D(key_mem_new[56]), .Z(key_mem_0__127__N_6112[56])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i57_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i60_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [59]), 
         .D(key_mem_new[59]), .Z(key_mem_0__127__N_6112[59])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i60_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i59_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [58]), 
         .D(key_mem_new[58]), .Z(key_mem_0__127__N_6112[58])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i59_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i62_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [61]), 
         .D(key_mem_new[61]), .Z(key_mem_0__127__N_6112[61])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i62_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i61_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [60]), 
         .D(key_mem_new[60]), .Z(key_mem_0__127__N_6112[60])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i61_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i10427 (.BLUT(n16017), .ALUT(n16022), .C0(n35835), .Z(n16023));
    LUT4 mux_14_i64_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [63]), 
         .D(key_mem_new[63]), .Z(key_mem_0__127__N_6112[63])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i64_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i63_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [62]), 
         .D(key_mem_new[62]), .Z(key_mem_0__127__N_6112[62])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i63_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i10488 (.BLUT(n16077), .ALUT(n16082), .C0(n35835), .Z(n16083));
    PFUMX i25744 (.BLUT(n1_adj_9005), .ALUT(n2_adj_9002), .C0(\muxed_round_nr[1] ), 
          .Z(n30903));
    LUT4 mux_14_i2_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [1]), 
         .D(key_mem_new[1]), .Z(key_mem_0__127__N_6112[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i1_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [0]), 
         .D(key_mem_new[0]), .Z(key_mem_0__127__N_6112[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i4_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [3]), 
         .D(key_mem_new[3]), .Z(key_mem_0__127__N_6112[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i3_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [2]), 
         .D(key_mem_new[2]), .Z(key_mem_0__127__N_6112[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i6_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [5]), 
         .D(key_mem_new[5]), .Z(key_mem_0__127__N_6112[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i5_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [4]), 
         .D(key_mem_new[4]), .Z(key_mem_0__127__N_6112[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i5_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25142 (.BLUT(n1_adj_9014), .ALUT(n2_adj_9012), .C0(\muxed_round_nr[1] ), 
          .Z(n30301));
    LUT4 mux_14_i8_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [7]), 
         .D(key_mem_new[7]), .Z(key_mem_0__127__N_6112[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i7_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [6]), 
         .D(key_mem_new[6]), .Z(key_mem_0__127__N_6112[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i10_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [9]), 
         .D(key_mem_new[9]), .Z(key_mem_0__127__N_6112[9])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i10_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i9_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [8]), 
         .D(key_mem_new[8]), .Z(key_mem_0__127__N_6112[8])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i9_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i12_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [11]), 
         .D(key_mem_new[11]), .Z(key_mem_0__127__N_6112[11])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i12_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i10549 (.BLUT(n16137), .ALUT(n16142), .C0(n35835), .Z(n16143));
    PFUMX i25143 (.BLUT(n4_adj_9010), .ALUT(n5_adj_9009), .C0(\muxed_round_nr[1] ), 
          .Z(n30302));
    LUT4 mux_14_i11_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [10]), 
         .D(key_mem_new[10]), .Z(key_mem_0__127__N_6112[10])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i11_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i10610 (.BLUT(n16197), .ALUT(n16202), .C0(n35835), .Z(n16203));
    LUT4 mux_14_i14_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [13]), 
         .D(key_mem_new[13]), .Z(key_mem_0__127__N_6112[13])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i14_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25144 (.BLUT(n8_adj_9008), .ALUT(n9_adj_9006), .C0(\muxed_round_nr[1] ), 
          .Z(n30303));
    LUT4 mux_14_i13_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [12]), 
         .D(key_mem_new[12]), .Z(key_mem_0__127__N_6112[12])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i13_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i16_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [15]), 
         .D(key_mem_new[15]), .Z(key_mem_0__127__N_6112[15])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i16_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i15_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [14]), 
         .D(key_mem_new[14]), .Z(key_mem_0__127__N_6112[14])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i15_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i18_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [17]), 
         .D(key_mem_new[17]), .Z(key_mem_0__127__N_6112[17])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i18_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i17_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [16]), 
         .D(key_mem_new[16]), .Z(key_mem_0__127__N_6112[16])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i17_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i20_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [19]), 
         .D(key_mem_new[19]), .Z(key_mem_0__127__N_6112[19])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i20_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i19_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [18]), 
         .D(key_mem_new[18]), .Z(key_mem_0__127__N_6112[18])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i19_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i22_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [21]), 
         .D(key_mem_new[21]), .Z(key_mem_0__127__N_6112[21])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i22_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i21_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [20]), 
         .D(key_mem_new[20]), .Z(key_mem_0__127__N_6112[20])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i21_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i10671 (.BLUT(n16257), .ALUT(n16262), .C0(n35835), .Z(n16263));
    LUT4 mux_14_i24_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [23]), 
         .D(key_mem_new[23]), .Z(key_mem_0__127__N_6112[23])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i24_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i23_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [22]), 
         .D(key_mem_new[22]), .Z(key_mem_0__127__N_6112[22])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i23_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i10732 (.BLUT(n16317), .ALUT(n16322), .C0(n35835), .Z(n16323));
    PFUMX i25149 (.BLUT(n1_adj_8999), .ALUT(n2_adj_8998), .C0(\muxed_round_nr[1] ), 
          .Z(n30308));
    LUT4 mux_14_i26_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [25]), 
         .D(key_mem_new[25]), .Z(key_mem_0__127__N_6112[25])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i26_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25745 (.BLUT(n4_adj_8991), .ALUT(n5_adj_8986), .C0(\muxed_round_nr[1] ), 
          .Z(n30904));
    LUT4 mux_14_i25_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [24]), 
         .D(key_mem_new[24]), .Z(key_mem_0__127__N_6112[24])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i25_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i28_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [27]), 
         .D(key_mem_new[27]), .Z(key_mem_0__127__N_6112[27])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i28_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i27_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [26]), 
         .D(key_mem_new[26]), .Z(key_mem_0__127__N_6112[26])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i27_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i30_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [29]), 
         .D(key_mem_new[29]), .Z(key_mem_0__127__N_6112[29])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i30_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i29_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [28]), 
         .D(key_mem_new[28]), .Z(key_mem_0__127__N_6112[28])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i29_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i32_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [31]), 
         .D(key_mem_new[31]), .Z(key_mem_0__127__N_6112[31])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i32_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i31_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [30]), 
         .D(key_mem_new[30]), .Z(key_mem_0__127__N_6112[30])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i31_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i10793 (.BLUT(n16377), .ALUT(n16382), .C0(n35835), .Z(n16383));
    LUT4 mux_14_i34_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [33]), 
         .D(key_mem_new[33]), .Z(key_mem_0__127__N_6112[33])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i34_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i33_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [32]), 
         .D(key_mem_new[32]), .Z(key_mem_0__127__N_6112[32])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i33_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i36_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [35]), 
         .D(key_mem_new[35]), .Z(key_mem_0__127__N_6112[35])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i36_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i35_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [34]), 
         .D(key_mem_new[34]), .Z(key_mem_0__127__N_6112[34])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i35_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i37_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [36]), 
         .D(key_mem_new[36]), .Z(key_mem_0__127__N_6112[36])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i37_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i66_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [65]), 
         .D(key_mem_new[65]), .Z(key_mem_0__127__N_6112[65])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i66_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i67_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [66]), 
         .D(key_mem_new[66]), .Z(key_mem_0__127__N_6112[66])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i67_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i68_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [67]), 
         .D(key_mem_new[67]), .Z(key_mem_0__127__N_6112[67])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i68_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i69_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [68]), 
         .D(key_mem_new[68]), .Z(key_mem_0__127__N_6112[68])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i69_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i70_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [69]), 
         .D(key_mem_new[69]), .Z(key_mem_0__127__N_6112[69])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i70_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i71_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [70]), 
         .D(key_mem_new[70]), .Z(key_mem_0__127__N_6112[70])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i71_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i72_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [71]), 
         .D(key_mem_new[71]), .Z(key_mem_0__127__N_6112[71])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i72_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25150 (.BLUT(n4_adj_8997), .ALUT(n5_adj_8996), .C0(\muxed_round_nr[1] ), 
          .Z(n30309));
    LUT4 mux_14_i73_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [72]), 
         .D(key_mem_new[72]), .Z(key_mem_0__127__N_6112[72])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i73_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i10854 (.BLUT(n16437), .ALUT(n16442), .C0(n35835), .Z(n16443));
    LUT4 mux_14_i74_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [73]), 
         .D(key_mem_new[73]), .Z(key_mem_0__127__N_6112[73])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i74_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i10915 (.BLUT(n16497), .ALUT(n16502), .C0(n35835), .Z(n16503));
    PFUMX i25151 (.BLUT(n8_adj_8994), .ALUT(n9_adj_8992), .C0(\muxed_round_nr[1] ), 
          .Z(n30310));
    LUT4 mux_14_i75_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [74]), 
         .D(key_mem_new[74]), .Z(key_mem_0__127__N_6112[74])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i75_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i76_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [75]), 
         .D(key_mem_new[75]), .Z(key_mem_0__127__N_6112[75])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i76_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i77_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [76]), 
         .D(key_mem_new[76]), .Z(key_mem_0__127__N_6112[76])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i77_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i78_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [77]), 
         .D(key_mem_new[77]), .Z(key_mem_0__127__N_6112[77])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i78_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i79_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [78]), 
         .D(key_mem_new[78]), .Z(key_mem_0__127__N_6112[78])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i79_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i80_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [79]), 
         .D(key_mem_new[79]), .Z(key_mem_0__127__N_6112[79])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i80_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i81_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [80]), 
         .D(key_mem_new[80]), .Z(key_mem_0__127__N_6112[80])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i81_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i82_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [81]), 
         .D(key_mem_new[81]), .Z(key_mem_0__127__N_6112[81])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i82_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i83_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [82]), 
         .D(key_mem_new[82]), .Z(key_mem_0__127__N_6112[82])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i83_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i84_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [83]), 
         .D(key_mem_new[83]), .Z(key_mem_0__127__N_6112[83])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i84_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i85_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [84]), 
         .D(key_mem_new[84]), .Z(key_mem_0__127__N_6112[84])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i85_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i10976 (.BLUT(n16557), .ALUT(n16562), .C0(n35835), .Z(n16563));
    LUT4 mux_14_i86_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [85]), 
         .D(key_mem_new[85]), .Z(key_mem_0__127__N_6112[85])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i86_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i87_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [86]), 
         .D(key_mem_new[86]), .Z(key_mem_0__127__N_6112[86])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i87_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i88_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [87]), 
         .D(key_mem_new[87]), .Z(key_mem_0__127__N_6112[87])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i88_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i89_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [88]), 
         .D(key_mem_new[88]), .Z(key_mem_0__127__N_6112[88])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i89_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i90_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [89]), 
         .D(key_mem_new[89]), .Z(key_mem_0__127__N_6112[89])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i90_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i91_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [90]), 
         .D(key_mem_new[90]), .Z(key_mem_0__127__N_6112[90])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i91_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i92_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [91]), 
         .D(key_mem_new[91]), .Z(key_mem_0__127__N_6112[91])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i92_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i93_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [92]), 
         .D(key_mem_new[92]), .Z(key_mem_0__127__N_6112[92])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i93_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i94_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [93]), 
         .D(key_mem_new[93]), .Z(key_mem_0__127__N_6112[93])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i94_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i95_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [94]), 
         .D(key_mem_new[94]), .Z(key_mem_0__127__N_6112[94])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i95_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i96_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [95]), 
         .D(key_mem_new[95]), .Z(key_mem_0__127__N_6112[95])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i96_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i97_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [96]), 
         .D(key_mem_new[96]), .Z(key_mem_0__127__N_6112[96])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i97_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i98_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [97]), 
         .D(key_mem_new[97]), .Z(key_mem_0__127__N_6112[97])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i98_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i99_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [98]), 
         .D(key_mem_new[98]), .Z(key_mem_0__127__N_6112[98])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i99_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i100_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [99]), 
         .D(key_mem_new[99]), .Z(key_mem_0__127__N_6112[99])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i100_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i11037 (.BLUT(n16617), .ALUT(n16622), .C0(n35835), .Z(n16623));
    LUT4 mux_14_i101_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [100]), 
         .D(key_mem_new[100]), .Z(key_mem_0__127__N_6112[100])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i101_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i102_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [101]), 
         .D(key_mem_new[101]), .Z(key_mem_0__127__N_6112[101])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i102_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25156 (.BLUT(n1_adj_8987), .ALUT(n2_adj_8985), .C0(\muxed_round_nr[1] ), 
          .Z(n30315));
    PFUMX i11098 (.BLUT(n16677), .ALUT(n16682), .C0(n35835), .Z(n16683));
    PFUMX i25157 (.BLUT(n4_adj_8983), .ALUT(n5_adj_8982), .C0(\muxed_round_nr[1] ), 
          .Z(n30316));
    PFUMX i25746 (.BLUT(n8_adj_8977), .ALUT(n9_adj_8976), .C0(\muxed_round_nr[1] ), 
          .Z(n30905));
    LUT4 mux_14_i103_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [102]), 
         .D(key_mem_new[102]), .Z(key_mem_0__127__N_6112[102])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i103_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i11159 (.BLUT(n16737), .ALUT(n16742), .C0(n35835), .Z(n16743));
    LUT4 mux_14_i104_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [103]), 
         .D(key_mem_new[103]), .Z(key_mem_0__127__N_6112[103])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i104_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25158 (.BLUT(n8_adj_8981), .ALUT(n9_adj_8979), .C0(\muxed_round_nr[1] ), 
          .Z(n30317));
    LUT4 mux_14_i105_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [104]), 
         .D(key_mem_new[104]), .Z(key_mem_0__127__N_6112[104])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i105_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i106_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [105]), 
         .D(key_mem_new[105]), .Z(key_mem_0__127__N_6112[105])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i106_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i107_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [106]), 
         .D(key_mem_new[106]), .Z(key_mem_0__127__N_6112[106])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i107_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i108_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [107]), 
         .D(key_mem_new[107]), .Z(key_mem_0__127__N_6112[107])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i108_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i109_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [108]), 
         .D(key_mem_new[108]), .Z(key_mem_0__127__N_6112[108])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i109_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i110_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [109]), 
         .D(key_mem_new[109]), .Z(key_mem_0__127__N_6112[109])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i110_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i111_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [110]), 
         .D(key_mem_new[110]), .Z(key_mem_0__127__N_6112[110])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i111_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i112_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [111]), 
         .D(key_mem_new[111]), .Z(key_mem_0__127__N_6112[111])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i112_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i113_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [112]), 
         .D(key_mem_new[112]), .Z(key_mem_0__127__N_6112[112])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i113_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25163 (.BLUT(n1_adj_8975), .ALUT(n2_adj_8974), .C0(\muxed_round_nr[1] ), 
          .Z(n30322));
    PFUMX i25164 (.BLUT(n4_adj_8973), .ALUT(n5_adj_8972), .C0(\muxed_round_nr[1] ), 
          .Z(n30323));
    LUT4 mux_14_i114_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [113]), 
         .D(key_mem_new[113]), .Z(key_mem_0__127__N_6112[113])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i114_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25165 (.BLUT(n8_adj_8971), .ALUT(n9_adj_8970), .C0(\muxed_round_nr[1] ), 
          .Z(n30324));
    LUT4 mux_14_i115_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [114]), 
         .D(key_mem_new[114]), .Z(key_mem_0__127__N_6112[114])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i115_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i116_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [115]), 
         .D(key_mem_new[115]), .Z(key_mem_0__127__N_6112[115])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i116_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i117_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [116]), 
         .D(key_mem_new[116]), .Z(key_mem_0__127__N_6112[116])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i117_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i118_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [117]), 
         .D(key_mem_new[117]), .Z(key_mem_0__127__N_6112[117])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i118_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i119_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [118]), 
         .D(key_mem_new[118]), .Z(key_mem_0__127__N_6112[118])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i119_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i120_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [119]), 
         .D(key_mem_new[119]), .Z(key_mem_0__127__N_6112[119])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i120_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i121_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [120]), 
         .D(key_mem_new[120]), .Z(key_mem_0__127__N_6112[120])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i121_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i122_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [121]), 
         .D(key_mem_new[121]), .Z(key_mem_0__127__N_6112[121])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i122_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i123_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [122]), 
         .D(key_mem_new[122]), .Z(key_mem_0__127__N_6112[122])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i123_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i124_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [123]), 
         .D(key_mem_new[123]), .Z(key_mem_0__127__N_6112[123])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i124_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i125_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [124]), 
         .D(key_mem_new[124]), .Z(key_mem_0__127__N_6112[124])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i125_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i126_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [125]), 
         .D(key_mem_new[125]), .Z(key_mem_0__127__N_6112[125])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i126_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i127_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [126]), 
         .D(key_mem_new[126]), .Z(key_mem_0__127__N_6112[126])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i127_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_14_i128_3_lut_4_lut (.A(n33945), .B(n33937), .C(\key_mem[9] [127]), 
         .D(key_mem_new[127]), .Z(key_mem_0__127__N_6112[127])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_14_i128_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i65_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [64]), 
         .D(key_mem_new[64]), .Z(key_mem_0__127__N_6240[64])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i65_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i39_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [38]), 
         .D(key_mem_new[38]), .Z(key_mem_0__127__N_6240[38])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i39_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i40_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [39]), 
         .D(key_mem_new[39]), .Z(key_mem_0__127__N_6240[39])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i40_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i41_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [40]), 
         .D(key_mem_new[40]), .Z(key_mem_0__127__N_6240[40])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i41_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i42_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [41]), 
         .D(key_mem_new[41]), .Z(key_mem_0__127__N_6240[41])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i42_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i43_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [42]), 
         .D(key_mem_new[42]), .Z(key_mem_0__127__N_6240[42])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i43_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i44_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [43]), 
         .D(key_mem_new[43]), .Z(key_mem_0__127__N_6240[43])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i44_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i45_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [44]), 
         .D(key_mem_new[44]), .Z(key_mem_0__127__N_6240[44])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i45_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i46_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [45]), 
         .D(key_mem_new[45]), .Z(key_mem_0__127__N_6240[45])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i46_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25170 (.BLUT(n1_adj_8967), .ALUT(n2_adj_8966), .C0(\muxed_round_nr[1] ), 
          .Z(n30329));
    LUT4 mux_13_i47_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [46]), 
         .D(key_mem_new[46]), .Z(key_mem_0__127__N_6240[46])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i47_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25171 (.BLUT(n4_adj_8965), .ALUT(n5_adj_8964), .C0(\muxed_round_nr[1] ), 
          .Z(n30330));
    LUT4 mux_13_i48_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [47]), 
         .D(key_mem_new[47]), .Z(key_mem_0__127__N_6240[47])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i48_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25172 (.BLUT(n8_adj_8963), .ALUT(n9_adj_8962), .C0(\muxed_round_nr[1] ), 
          .Z(n30331));
    LUT4 mux_13_i49_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [48]), 
         .D(key_mem_new[48]), .Z(key_mem_0__127__N_6240[48])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i49_3_lut_4_lut.init = 16'hf1e0;
    PFUMX keylen_I_0_Mux_127_i1 (.BLUT(key_mem_new_127__N_7264[127]), .ALUT(prev_key1_new_127__N_7520[127]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[127])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    LUT4 mux_13_i50_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [49]), 
         .D(key_mem_new[49]), .Z(key_mem_0__127__N_6240[49])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i50_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i51_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [50]), 
         .D(key_mem_new[50]), .Z(key_mem_0__127__N_6240[50])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i51_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25177 (.BLUT(n1_adj_8960), .ALUT(n2_adj_8959), .C0(\muxed_round_nr[1] ), 
          .Z(n30336));
    PFUMX keylen_I_0_Mux_126_i1 (.BLUT(key_mem_new_127__N_7264[126]), .ALUT(prev_key1_new_127__N_7520[126]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[126])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    LUT4 mux_13_i52_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [51]), 
         .D(key_mem_new[51]), .Z(key_mem_0__127__N_6240[51])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i52_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i53_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [52]), 
         .D(key_mem_new[52]), .Z(key_mem_0__127__N_6240[52])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i53_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i54_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [53]), 
         .D(key_mem_new[53]), .Z(key_mem_0__127__N_6240[53])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i54_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i55_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [54]), 
         .D(key_mem_new[54]), .Z(key_mem_0__127__N_6240[54])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i55_3_lut_4_lut.init = 16'hf1e0;
    PFUMX keylen_I_0_Mux_125_i1 (.BLUT(key_mem_new_127__N_7264[125]), .ALUT(prev_key1_new_127__N_7520[125]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[125])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    PFUMX i25751 (.BLUT(n1_adj_8958), .ALUT(n2_adj_8955), .C0(\muxed_round_nr[1] ), 
          .Z(n30910));
    LUT4 mux_13_i56_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [55]), 
         .D(key_mem_new[55]), .Z(key_mem_0__127__N_6240[55])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i56_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i57_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [56]), 
         .D(key_mem_new[56]), .Z(key_mem_0__127__N_6240[56])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i57_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i58_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [57]), 
         .D(key_mem_new[57]), .Z(key_mem_0__127__N_6240[57])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i58_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i59_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [58]), 
         .D(key_mem_new[58]), .Z(key_mem_0__127__N_6240[58])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i59_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i60_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [59]), 
         .D(key_mem_new[59]), .Z(key_mem_0__127__N_6240[59])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i60_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i61_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [60]), 
         .D(key_mem_new[60]), .Z(key_mem_0__127__N_6240[60])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i61_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25178 (.BLUT(n4_adj_8954), .ALUT(n5_adj_8951), .C0(\muxed_round_nr[1] ), 
          .Z(n30337));
    LUT4 mux_13_i62_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [61]), 
         .D(key_mem_new[61]), .Z(key_mem_0__127__N_6240[61])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i62_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i63_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [62]), 
         .D(key_mem_new[62]), .Z(key_mem_0__127__N_6240[62])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i63_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i64_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [63]), 
         .D(key_mem_new[63]), .Z(key_mem_0__127__N_6240[63])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i64_3_lut_4_lut.init = 16'hf1e0;
    PFUMX keylen_I_0_Mux_124_i1 (.BLUT(key_mem_new_127__N_7264[124]), .ALUT(prev_key1_new_127__N_7520[124]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[124])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    LUT4 mux_13_i1_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [0]), 
         .D(key_mem_new[0]), .Z(key_mem_0__127__N_6240[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i2_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [1]), 
         .D(key_mem_new[1]), .Z(key_mem_0__127__N_6240[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i3_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [2]), 
         .D(key_mem_new[2]), .Z(key_mem_0__127__N_6240[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i4_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [3]), 
         .D(key_mem_new[3]), .Z(key_mem_0__127__N_6240[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i5_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [4]), 
         .D(key_mem_new[4]), .Z(key_mem_0__127__N_6240[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i6_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [5]), 
         .D(key_mem_new[5]), .Z(key_mem_0__127__N_6240[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i7_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [6]), 
         .D(key_mem_new[6]), .Z(key_mem_0__127__N_6240[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i8_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [7]), 
         .D(key_mem_new[7]), .Z(key_mem_0__127__N_6240[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i8_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25752 (.BLUT(n4_adj_8953), .ALUT(n5_adj_8952), .C0(\muxed_round_nr[1] ), 
          .Z(n30911));
    PFUMX keylen_I_0_Mux_123_i1 (.BLUT(key_mem_new_127__N_7264[123]), .ALUT(prev_key1_new_127__N_7520[123]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[123])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    LUT4 mux_13_i9_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [8]), 
         .D(key_mem_new[8]), .Z(key_mem_0__127__N_6240[8])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i9_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i10_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [9]), 
         .D(key_mem_new[9]), .Z(key_mem_0__127__N_6240[9])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i10_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i11_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [10]), 
         .D(key_mem_new[10]), .Z(key_mem_0__127__N_6240[10])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i11_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i12_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [11]), 
         .D(key_mem_new[11]), .Z(key_mem_0__127__N_6240[11])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i12_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25179 (.BLUT(n8_adj_8950), .ALUT(n9_adj_8949), .C0(\muxed_round_nr[1] ), 
          .Z(n30338));
    LUT4 mux_13_i13_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [12]), 
         .D(key_mem_new[12]), .Z(key_mem_0__127__N_6240[12])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i13_3_lut_4_lut.init = 16'hf1e0;
    PFUMX keylen_I_0_Mux_122_i1 (.BLUT(key_mem_new_127__N_7264[122]), .ALUT(prev_key1_new_127__N_7520[122]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[122])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    LUT4 mux_13_i14_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [13]), 
         .D(key_mem_new[13]), .Z(key_mem_0__127__N_6240[13])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i14_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i15_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [14]), 
         .D(key_mem_new[14]), .Z(key_mem_0__127__N_6240[14])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i15_3_lut_4_lut.init = 16'hf1e0;
    PFUMX keylen_I_0_Mux_121_i1 (.BLUT(key_mem_new_127__N_7264[121]), .ALUT(prev_key1_new_127__N_7520[121]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[121])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    LUT4 mux_13_i16_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [15]), 
         .D(key_mem_new[15]), .Z(key_mem_0__127__N_6240[15])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i16_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i17_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [16]), 
         .D(key_mem_new[16]), .Z(key_mem_0__127__N_6240[16])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i17_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25753 (.BLUT(n8_adj_8947), .ALUT(n9_adj_8941), .C0(\muxed_round_nr[1] ), 
          .Z(n30912));
    LUT4 mux_13_i18_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [17]), 
         .D(key_mem_new[17]), .Z(key_mem_0__127__N_6240[17])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i18_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i19_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [18]), 
         .D(key_mem_new[18]), .Z(key_mem_0__127__N_6240[18])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i19_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i20_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [19]), 
         .D(key_mem_new[19]), .Z(key_mem_0__127__N_6240[19])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i20_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25184 (.BLUT(n1_adj_8946), .ALUT(n2_adj_8945), .C0(\muxed_round_nr[1] ), 
          .Z(n30343));
    PFUMX keylen_I_0_Mux_120_i1 (.BLUT(key_mem_new_127__N_7264[120]), .ALUT(prev_key1_new_127__N_7520[120]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[120])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    LUT4 mux_13_i21_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [20]), 
         .D(key_mem_new[20]), .Z(key_mem_0__127__N_6240[20])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i21_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25185 (.BLUT(n4_adj_8944), .ALUT(n5_adj_8943), .C0(\muxed_round_nr[1] ), 
          .Z(n30344));
    LUT4 mux_13_i22_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [21]), 
         .D(key_mem_new[21]), .Z(key_mem_0__127__N_6240[21])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i22_3_lut_4_lut.init = 16'hf1e0;
    PFUMX keylen_I_0_Mux_87_i1 (.BLUT(key_mem_new_127__N_7264[87]), .ALUT(prev_key1_new_127__N_7520[87]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[87])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    LUT4 mux_13_i23_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [22]), 
         .D(key_mem_new[22]), .Z(key_mem_0__127__N_6240[22])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i23_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i24_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [23]), 
         .D(key_mem_new[23]), .Z(key_mem_0__127__N_6240[23])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i24_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i25_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [24]), 
         .D(key_mem_new[24]), .Z(key_mem_0__127__N_6240[24])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i25_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i26_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [25]), 
         .D(key_mem_new[25]), .Z(key_mem_0__127__N_6240[25])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i26_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i27_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [26]), 
         .D(key_mem_new[26]), .Z(key_mem_0__127__N_6240[26])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i27_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i28_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [27]), 
         .D(key_mem_new[27]), .Z(key_mem_0__127__N_6240[27])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i28_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i29_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [28]), 
         .D(key_mem_new[28]), .Z(key_mem_0__127__N_6240[28])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i29_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i30_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [29]), 
         .D(key_mem_new[29]), .Z(key_mem_0__127__N_6240[29])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i30_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i31_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [30]), 
         .D(key_mem_new[30]), .Z(key_mem_0__127__N_6240[30])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i31_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i32_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [31]), 
         .D(key_mem_new[31]), .Z(key_mem_0__127__N_6240[31])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i32_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i33_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [32]), 
         .D(key_mem_new[32]), .Z(key_mem_0__127__N_6240[32])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i33_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i34_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [33]), 
         .D(key_mem_new[33]), .Z(key_mem_0__127__N_6240[33])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i34_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25186 (.BLUT(n8_adj_8942), .ALUT(n9_adj_8940), .C0(\muxed_round_nr[1] ), 
          .Z(n30345));
    LUT4 mux_13_i35_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [34]), 
         .D(key_mem_new[34]), .Z(key_mem_0__127__N_6240[34])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i35_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i36_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [35]), 
         .D(key_mem_new[35]), .Z(key_mem_0__127__N_6240[35])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i36_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i37_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [36]), 
         .D(key_mem_new[36]), .Z(key_mem_0__127__N_6240[36])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i37_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i38_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [37]), 
         .D(key_mem_new[37]), .Z(key_mem_0__127__N_6240[37])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i38_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i66_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [65]), 
         .D(key_mem_new[65]), .Z(key_mem_0__127__N_6240[65])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i66_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i67_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [66]), 
         .D(key_mem_new[66]), .Z(key_mem_0__127__N_6240[66])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i67_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i68_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [67]), 
         .D(key_mem_new[67]), .Z(key_mem_0__127__N_6240[67])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i68_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i69_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [68]), 
         .D(key_mem_new[68]), .Z(key_mem_0__127__N_6240[68])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i69_3_lut_4_lut.init = 16'hf1e0;
    PFUMX keylen_I_0_Mux_86_i1 (.BLUT(key_mem_new_127__N_7264[86]), .ALUT(prev_key1_new_127__N_7520[86]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[86])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    LUT4 mux_13_i70_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [69]), 
         .D(key_mem_new[69]), .Z(key_mem_0__127__N_6240[69])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i70_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i71_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [70]), 
         .D(key_mem_new[70]), .Z(key_mem_0__127__N_6240[70])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i71_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25191 (.BLUT(n1_adj_8938), .ALUT(n2_adj_8937), .C0(\muxed_round_nr[1] ), 
          .Z(n30350));
    PFUMX keylen_I_0_Mux_85_i1 (.BLUT(key_mem_new_127__N_7264[85]), .ALUT(prev_key1_new_127__N_7520[85]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[85])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    LUT4 mux_13_i72_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [71]), 
         .D(key_mem_new[71]), .Z(key_mem_0__127__N_6240[71])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i72_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i73_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [72]), 
         .D(key_mem_new[72]), .Z(key_mem_0__127__N_6240[72])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i73_3_lut_4_lut.init = 16'hf1e0;
    PFUMX keylen_I_0_Mux_84_i1 (.BLUT(key_mem_new_127__N_7264[84]), .ALUT(prev_key1_new_127__N_7520[84]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[84])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    PFUMX i25192 (.BLUT(n4_adj_8936), .ALUT(n5_adj_8934), .C0(\muxed_round_nr[1] ), 
          .Z(n30351));
    LUT4 mux_13_i74_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [73]), 
         .D(key_mem_new[73]), .Z(key_mem_0__127__N_6240[73])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i74_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i75_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [74]), 
         .D(key_mem_new[74]), .Z(key_mem_0__127__N_6240[74])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i75_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i76_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [75]), 
         .D(key_mem_new[75]), .Z(key_mem_0__127__N_6240[75])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i76_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i77_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [76]), 
         .D(key_mem_new[76]), .Z(key_mem_0__127__N_6240[76])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i77_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25193 (.BLUT(n8_adj_8933), .ALUT(n9_adj_8932), .C0(\muxed_round_nr[1] ), 
          .Z(n30352));
    LUT4 mux_13_i78_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [77]), 
         .D(key_mem_new[77]), .Z(key_mem_0__127__N_6240[77])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i78_3_lut_4_lut.init = 16'hf1e0;
    PFUMX keylen_I_0_Mux_83_i1 (.BLUT(key_mem_new_127__N_7264[83]), .ALUT(prev_key1_new_127__N_7520[83]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[83])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    LUT4 mux_13_i79_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [78]), 
         .D(key_mem_new[78]), .Z(key_mem_0__127__N_6240[78])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i79_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i80_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [79]), 
         .D(key_mem_new[79]), .Z(key_mem_0__127__N_6240[79])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i80_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25758 (.BLUT(n1_adj_8931), .ALUT(n2_adj_8930), .C0(\muxed_round_nr[1] ), 
          .Z(n30917));
    LUT4 mux_13_i81_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [80]), 
         .D(key_mem_new[80]), .Z(key_mem_0__127__N_6240[80])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i81_3_lut_4_lut.init = 16'hf1e0;
    PFUMX keylen_I_0_Mux_82_i1 (.BLUT(key_mem_new_127__N_7264[82]), .ALUT(prev_key1_new_127__N_7520[82]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[82])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    LUT4 mux_13_i82_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [81]), 
         .D(key_mem_new[81]), .Z(key_mem_0__127__N_6240[81])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i82_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i83_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [82]), 
         .D(key_mem_new[82]), .Z(key_mem_0__127__N_6240[82])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i83_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i84_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [83]), 
         .D(key_mem_new[83]), .Z(key_mem_0__127__N_6240[83])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i84_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i85_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [84]), 
         .D(key_mem_new[84]), .Z(key_mem_0__127__N_6240[84])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i85_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i86_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [85]), 
         .D(key_mem_new[85]), .Z(key_mem_0__127__N_6240[85])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i86_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i87_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [86]), 
         .D(key_mem_new[86]), .Z(key_mem_0__127__N_6240[86])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i87_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i88_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [87]), 
         .D(key_mem_new[87]), .Z(key_mem_0__127__N_6240[87])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i88_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i89_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [88]), 
         .D(key_mem_new[88]), .Z(key_mem_0__127__N_6240[88])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i89_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i90_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [89]), 
         .D(key_mem_new[89]), .Z(key_mem_0__127__N_6240[89])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i90_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i91_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [90]), 
         .D(key_mem_new[90]), .Z(key_mem_0__127__N_6240[90])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i91_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i92_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [91]), 
         .D(key_mem_new[91]), .Z(key_mem_0__127__N_6240[91])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i92_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i93_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [92]), 
         .D(key_mem_new[92]), .Z(key_mem_0__127__N_6240[92])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i93_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i94_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [93]), 
         .D(key_mem_new[93]), .Z(key_mem_0__127__N_6240[93])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i94_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i95_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [94]), 
         .D(key_mem_new[94]), .Z(key_mem_0__127__N_6240[94])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i95_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i96_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [95]), 
         .D(key_mem_new[95]), .Z(key_mem_0__127__N_6240[95])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i96_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i97_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [96]), 
         .D(key_mem_new[96]), .Z(key_mem_0__127__N_6240[96])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i97_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i98_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [97]), 
         .D(key_mem_new[97]), .Z(key_mem_0__127__N_6240[97])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i98_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i99_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [98]), 
         .D(key_mem_new[98]), .Z(key_mem_0__127__N_6240[98])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i99_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i100_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [99]), 
         .D(key_mem_new[99]), .Z(key_mem_0__127__N_6240[99])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i100_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i101_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [100]), 
         .D(key_mem_new[100]), .Z(key_mem_0__127__N_6240[100])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i101_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i102_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [101]), 
         .D(key_mem_new[101]), .Z(key_mem_0__127__N_6240[101])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i102_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i103_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [102]), 
         .D(key_mem_new[102]), .Z(key_mem_0__127__N_6240[102])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i103_3_lut_4_lut.init = 16'hf1e0;
    PFUMX keylen_I_0_Mux_81_i1 (.BLUT(key_mem_new_127__N_7264[81]), .ALUT(prev_key1_new_127__N_7520[81]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[81])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    LUT4 mux_13_i104_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [103]), 
         .D(key_mem_new[103]), .Z(key_mem_0__127__N_6240[103])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i104_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i105_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [104]), 
         .D(key_mem_new[104]), .Z(key_mem_0__127__N_6240[104])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i105_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i106_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [105]), 
         .D(key_mem_new[105]), .Z(key_mem_0__127__N_6240[105])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i106_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i107_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [106]), 
         .D(key_mem_new[106]), .Z(key_mem_0__127__N_6240[106])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i107_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i108_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [107]), 
         .D(key_mem_new[107]), .Z(key_mem_0__127__N_6240[107])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i108_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i109_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [108]), 
         .D(key_mem_new[108]), .Z(key_mem_0__127__N_6240[108])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i109_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i110_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [109]), 
         .D(key_mem_new[109]), .Z(key_mem_0__127__N_6240[109])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i110_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i111_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [110]), 
         .D(key_mem_new[110]), .Z(key_mem_0__127__N_6240[110])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i111_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i112_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [111]), 
         .D(key_mem_new[111]), .Z(key_mem_0__127__N_6240[111])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i112_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i113_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [112]), 
         .D(key_mem_new[112]), .Z(key_mem_0__127__N_6240[112])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i113_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i114_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [113]), 
         .D(key_mem_new[113]), .Z(key_mem_0__127__N_6240[113])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i114_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i115_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [114]), 
         .D(key_mem_new[114]), .Z(key_mem_0__127__N_6240[114])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i115_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i116_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [115]), 
         .D(key_mem_new[115]), .Z(key_mem_0__127__N_6240[115])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i116_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i117_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [116]), 
         .D(key_mem_new[116]), .Z(key_mem_0__127__N_6240[116])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i117_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i118_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [117]), 
         .D(key_mem_new[117]), .Z(key_mem_0__127__N_6240[117])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i118_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i119_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [118]), 
         .D(key_mem_new[118]), .Z(key_mem_0__127__N_6240[118])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i119_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i120_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [119]), 
         .D(key_mem_new[119]), .Z(key_mem_0__127__N_6240[119])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i120_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i121_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [120]), 
         .D(key_mem_new[120]), .Z(key_mem_0__127__N_6240[120])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i121_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i122_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [121]), 
         .D(key_mem_new[121]), .Z(key_mem_0__127__N_6240[121])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i122_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i123_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [122]), 
         .D(key_mem_new[122]), .Z(key_mem_0__127__N_6240[122])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i123_3_lut_4_lut.init = 16'hf1e0;
    PFUMX keylen_I_0_Mux_80_i1 (.BLUT(key_mem_new_127__N_7264[80]), .ALUT(prev_key1_new_127__N_7520[80]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[80])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    LUT4 mux_13_i124_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [123]), 
         .D(key_mem_new[123]), .Z(key_mem_0__127__N_6240[123])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i124_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i125_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [124]), 
         .D(key_mem_new[124]), .Z(key_mem_0__127__N_6240[124])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i125_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i126_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [125]), 
         .D(key_mem_new[125]), .Z(key_mem_0__127__N_6240[125])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i126_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_13_i127_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [126]), 
         .D(key_mem_new[126]), .Z(key_mem_0__127__N_6240[126])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i127_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25759 (.BLUT(n4_adj_8928), .ALUT(n5_adj_8927), .C0(\muxed_round_nr[1] ), 
          .Z(n30918));
    PFUMX i25198 (.BLUT(n1_adj_8926), .ALUT(n2_adj_8925), .C0(\muxed_round_nr[1] ), 
          .Z(n30357));
    LUT4 mux_13_i128_3_lut_4_lut (.A(n33912), .B(n33937), .C(\key_mem[10] [127]), 
         .D(key_mem_new[127]), .Z(key_mem_0__127__N_6240[127])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_13_i128_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_12_i65_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [64]), 
         .D(key_mem_new[64]), .Z(key_mem_0__127__N_6368[64])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i65_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25760 (.BLUT(n8_adj_8924), .ALUT(n9_adj_8923), .C0(\muxed_round_nr[1] ), 
          .Z(n30919));
    PFUMX keylen_I_0_Mux_79_i1 (.BLUT(key_mem_new_127__N_7264[79]), .ALUT(prev_key1_new_127__N_7520[79]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[79])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    LUT4 mux_12_i40_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [39]), 
         .D(key_mem_new[39]), .Z(key_mem_0__127__N_6368[39])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i40_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25199 (.BLUT(n4_adj_8922), .ALUT(n5_adj_8920), .C0(\muxed_round_nr[1] ), 
          .Z(n30358));
    LUT4 mux_12_i41_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [40]), 
         .D(key_mem_new[40]), .Z(key_mem_0__127__N_6368[40])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i41_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i42_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [41]), 
         .D(key_mem_new[41]), .Z(key_mem_0__127__N_6368[41])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i42_3_lut_4_lut.init = 16'hf2d0;
    PFUMX keylen_I_0_Mux_78_i1 (.BLUT(key_mem_new_127__N_7264[78]), .ALUT(prev_key1_new_127__N_7520[78]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[78])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    PFUMX i25862 (.BLUT(n4_adj_8919), .ALUT(n5_adj_8918), .C0(\muxed_round_nr[1] ), 
          .Z(n31021));
    PFUMX i25200 (.BLUT(n8_adj_8916), .ALUT(n9_adj_8914), .C0(\muxed_round_nr[1] ), 
          .Z(n30359));
    LUT4 mux_12_i43_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [42]), 
         .D(key_mem_new[42]), .Z(key_mem_0__127__N_6368[42])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i43_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i44_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [43]), 
         .D(key_mem_new[43]), .Z(key_mem_0__127__N_6368[43])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i44_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i45_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [44]), 
         .D(key_mem_new[44]), .Z(key_mem_0__127__N_6368[44])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i45_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i46_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [45]), 
         .D(key_mem_new[45]), .Z(key_mem_0__127__N_6368[45])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i46_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25863 (.BLUT(n8_adj_8917), .ALUT(n9_adj_8915), .C0(\muxed_round_nr[1] ), 
          .Z(n31022));
    LUT4 mux_12_i47_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [46]), 
         .D(key_mem_new[46]), .Z(key_mem_0__127__N_6368[46])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i47_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i48_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [47]), 
         .D(key_mem_new[47]), .Z(key_mem_0__127__N_6368[47])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i48_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i49_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [48]), 
         .D(key_mem_new[48]), .Z(key_mem_0__127__N_6368[48])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i49_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i50_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [49]), 
         .D(key_mem_new[49]), .Z(key_mem_0__127__N_6368[49])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i50_3_lut_4_lut.init = 16'hf2d0;
    PFUMX keylen_I_0_Mux_77_i1 (.BLUT(key_mem_new_127__N_7264[77]), .ALUT(prev_key1_new_127__N_7520[77]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[77])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    LUT4 mux_12_i51_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [50]), 
         .D(key_mem_new[50]), .Z(key_mem_0__127__N_6368[50])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i51_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i52_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [51]), 
         .D(key_mem_new[51]), .Z(key_mem_0__127__N_6368[51])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i52_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i53_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [52]), 
         .D(key_mem_new[52]), .Z(key_mem_0__127__N_6368[52])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i53_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25868 (.BLUT(n1_adj_8911), .ALUT(n2_adj_8910), .C0(\muxed_round_nr[1] ), 
          .Z(n31027));
    PFUMX keylen_I_0_Mux_76_i1 (.BLUT(key_mem_new_127__N_7264[76]), .ALUT(prev_key1_new_127__N_7520[76]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[76])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    PFUMX i25869 (.BLUT(n4_adj_8909), .ALUT(n5_adj_8908), .C0(\muxed_round_nr[1] ), 
          .Z(n31028));
    LUT4 mux_12_i54_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [53]), 
         .D(key_mem_new[53]), .Z(key_mem_0__127__N_6368[53])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i54_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i55_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [54]), 
         .D(key_mem_new[54]), .Z(key_mem_0__127__N_6368[54])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i55_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i56_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [55]), 
         .D(key_mem_new[55]), .Z(key_mem_0__127__N_6368[55])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i56_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25205 (.BLUT(n1_adj_8907), .ALUT(n2_adj_8905), .C0(\muxed_round_nr[1] ), 
          .Z(n30364));
    PFUMX keylen_I_0_Mux_75_i1 (.BLUT(key_mem_new_127__N_7264[75]), .ALUT(prev_key1_new_127__N_7520[75]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[75])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    PFUMX i25870 (.BLUT(n8_adj_8906), .ALUT(n9_adj_8904), .C0(\muxed_round_nr[1] ), 
          .Z(n31029));
    LUT4 mux_12_i57_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [56]), 
         .D(key_mem_new[56]), .Z(key_mem_0__127__N_6368[56])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i57_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i58_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [57]), 
         .D(key_mem_new[57]), .Z(key_mem_0__127__N_6368[57])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i58_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25206 (.BLUT(n4_adj_8903), .ALUT(n5_adj_8902), .C0(\muxed_round_nr[1] ), 
          .Z(n30365));
    LUT4 mux_12_i59_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [58]), 
         .D(key_mem_new[58]), .Z(key_mem_0__127__N_6368[58])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i59_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i60_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [59]), 
         .D(key_mem_new[59]), .Z(key_mem_0__127__N_6368[59])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i60_3_lut_4_lut.init = 16'hf2d0;
    PFUMX keylen_I_0_Mux_74_i1 (.BLUT(key_mem_new_127__N_7264[74]), .ALUT(prev_key1_new_127__N_7520[74]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[74])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    LUT4 mux_12_i61_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [60]), 
         .D(key_mem_new[60]), .Z(key_mem_0__127__N_6368[60])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i61_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i62_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [61]), 
         .D(key_mem_new[61]), .Z(key_mem_0__127__N_6368[61])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i62_3_lut_4_lut.init = 16'hf2d0;
    PFUMX keylen_I_0_Mux_73_i1 (.BLUT(key_mem_new_127__N_7264[73]), .ALUT(prev_key1_new_127__N_7520[73]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[73])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    PFUMX i25207 (.BLUT(n8_adj_8900), .ALUT(n9_adj_8898), .C0(\muxed_round_nr[1] ), 
          .Z(n30366));
    LUT4 mux_12_i63_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [62]), 
         .D(key_mem_new[62]), .Z(key_mem_0__127__N_6368[62])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i63_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25875 (.BLUT(n1_adj_8899), .ALUT(n2_adj_8897), .C0(\muxed_round_nr[1] ), 
          .Z(n31034));
    LUT4 mux_12_i64_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [63]), 
         .D(key_mem_new[63]), .Z(key_mem_0__127__N_6368[63])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i64_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i1_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [0]), 
         .D(key_mem_new[0]), .Z(key_mem_0__127__N_6368[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i1_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i2_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [1]), 
         .D(key_mem_new[1]), .Z(key_mem_0__127__N_6368[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i2_3_lut_4_lut.init = 16'hf2d0;
    PFUMX keylen_I_0_Mux_72_i1 (.BLUT(key_mem_new_127__N_7264[72]), .ALUT(prev_key1_new_127__N_7520[72]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[72])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    LUT4 mux_12_i3_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [2]), 
         .D(key_mem_new[2]), .Z(key_mem_0__127__N_6368[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i3_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i4_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [3]), 
         .D(key_mem_new[3]), .Z(key_mem_0__127__N_6368[3])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i4_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i5_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [4]), 
         .D(key_mem_new[4]), .Z(key_mem_0__127__N_6368[4])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i5_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i6_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [5]), 
         .D(key_mem_new[5]), .Z(key_mem_0__127__N_6368[5])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i6_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i7_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [6]), 
         .D(key_mem_new[6]), .Z(key_mem_0__127__N_6368[6])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i7_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i8_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [7]), 
         .D(key_mem_new[7]), .Z(key_mem_0__127__N_6368[7])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i8_3_lut_4_lut.init = 16'hf2d0;
    PFUMX keylen_I_0_Mux_71_i1 (.BLUT(key_mem_new_127__N_7264[71]), .ALUT(prev_key1_new_127__N_7520[71]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[71])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    LUT4 mux_12_i9_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [8]), 
         .D(key_mem_new[8]), .Z(key_mem_0__127__N_6368[8])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i9_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i10_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [9]), 
         .D(key_mem_new[9]), .Z(key_mem_0__127__N_6368[9])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i10_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25876 (.BLUT(n4_adj_8895), .ALUT(n5_adj_8894), .C0(\muxed_round_nr[1] ), 
          .Z(n31035));
    LUT4 mux_12_i11_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [10]), 
         .D(key_mem_new[10]), .Z(key_mem_0__127__N_6368[10])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i11_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i12_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [11]), 
         .D(key_mem_new[11]), .Z(key_mem_0__127__N_6368[11])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i12_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25212 (.BLUT(n1_adj_8893), .ALUT(n2_adj_8891), .C0(\muxed_round_nr[1] ), 
          .Z(n30371));
    PFUMX i25877 (.BLUT(n8_adj_8892), .ALUT(n9_adj_8890), .C0(\muxed_round_nr[1] ), 
          .Z(n31036));
    PFUMX keylen_I_0_Mux_70_i1 (.BLUT(key_mem_new_127__N_7264[70]), .ALUT(prev_key1_new_127__N_7520[70]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[70])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    LUT4 mux_12_i13_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [12]), 
         .D(key_mem_new[12]), .Z(key_mem_0__127__N_6368[12])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i13_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25213 (.BLUT(n4_adj_8889), .ALUT(n5_adj_8888), .C0(\muxed_round_nr[1] ), 
          .Z(n30372));
    LUT4 mux_12_i14_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [13]), 
         .D(key_mem_new[13]), .Z(key_mem_0__127__N_6368[13])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i14_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i15_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [14]), 
         .D(key_mem_new[14]), .Z(key_mem_0__127__N_6368[14])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i15_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i16_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [15]), 
         .D(key_mem_new[15]), .Z(key_mem_0__127__N_6368[15])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i16_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i17_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [16]), 
         .D(key_mem_new[16]), .Z(key_mem_0__127__N_6368[16])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i17_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i18_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [17]), 
         .D(key_mem_new[17]), .Z(key_mem_0__127__N_6368[17])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i18_3_lut_4_lut.init = 16'hf2d0;
    PFUMX keylen_I_0_Mux_69_i1 (.BLUT(key_mem_new_127__N_7264[69]), .ALUT(prev_key1_new_127__N_7520[69]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[69])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    PFUMX i25214 (.BLUT(n8_adj_8886), .ALUT(n9_adj_8883), .C0(\muxed_round_nr[1] ), 
          .Z(n30373));
    PFUMX i25882 (.BLUT(n1_adj_8885), .ALUT(n2_adj_8884), .C0(\muxed_round_nr[1] ), 
          .Z(n31041));
    LUT4 mux_12_i19_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [18]), 
         .D(key_mem_new[18]), .Z(key_mem_0__127__N_6368[18])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i19_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i20_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [19]), 
         .D(key_mem_new[19]), .Z(key_mem_0__127__N_6368[19])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i20_3_lut_4_lut.init = 16'hf2d0;
    PFUMX keylen_I_0_Mux_68_i1 (.BLUT(key_mem_new_127__N_7264[68]), .ALUT(prev_key1_new_127__N_7520[68]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[68])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    PFUMX i25883 (.BLUT(n4_adj_8882), .ALUT(n5_adj_8881), .C0(\muxed_round_nr[1] ), 
          .Z(n31042));
    LUT4 mux_12_i21_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [20]), 
         .D(key_mem_new[20]), .Z(key_mem_0__127__N_6368[20])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i21_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i22_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [21]), 
         .D(key_mem_new[21]), .Z(key_mem_0__127__N_6368[21])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i22_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i23_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [22]), 
         .D(key_mem_new[22]), .Z(key_mem_0__127__N_6368[22])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i23_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25884 (.BLUT(n8_adj_8879), .ALUT(n9_adj_8878), .C0(\muxed_round_nr[1] ), 
          .Z(n31043));
    PFUMX keylen_I_0_Mux_67_i1 (.BLUT(key_mem_new_127__N_7264[67]), .ALUT(prev_key1_new_127__N_7520[67]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[67])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    LUT4 mux_12_i24_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [23]), 
         .D(key_mem_new[23]), .Z(key_mem_0__127__N_6368[23])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i24_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i25_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [24]), 
         .D(key_mem_new[24]), .Z(key_mem_0__127__N_6368[24])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i25_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25219 (.BLUT(n1_adj_8876), .ALUT(n2_adj_8875), .C0(\muxed_round_nr[1] ), 
          .Z(n30378));
    LUT4 mux_12_i26_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [25]), 
         .D(key_mem_new[25]), .Z(key_mem_0__127__N_6368[25])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i26_3_lut_4_lut.init = 16'hf2d0;
    PFUMX keylen_I_0_Mux_66_i1 (.BLUT(key_mem_new_127__N_7264[66]), .ALUT(prev_key1_new_127__N_7520[66]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[66])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    PFUMX i25889 (.BLUT(n1_adj_8874), .ALUT(n2_adj_8873), .C0(\muxed_round_nr[1] ), 
          .Z(n31048));
    LUT4 mux_12_i27_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [26]), 
         .D(key_mem_new[26]), .Z(key_mem_0__127__N_6368[26])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i27_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i28_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [27]), 
         .D(key_mem_new[27]), .Z(key_mem_0__127__N_6368[27])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i28_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25220 (.BLUT(n4_adj_8872), .ALUT(n5_adj_8869), .C0(\muxed_round_nr[1] ), 
          .Z(n30379));
    PFUMX i25890 (.BLUT(n4_adj_8871), .ALUT(n5_adj_8870), .C0(\muxed_round_nr[1] ), 
          .Z(n31049));
    LUT4 mux_12_i29_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [28]), 
         .D(key_mem_new[28]), .Z(key_mem_0__127__N_6368[28])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i29_3_lut_4_lut.init = 16'hf2d0;
    PFUMX keylen_I_0_Mux_65_i1 (.BLUT(key_mem_new_127__N_7264[65]), .ALUT(prev_key1_new_127__N_7520[65]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[65])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    LUT4 mux_12_i30_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [29]), 
         .D(key_mem_new[29]), .Z(key_mem_0__127__N_6368[29])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i30_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i31_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [30]), 
         .D(key_mem_new[30]), .Z(key_mem_0__127__N_6368[30])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i31_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i32_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [31]), 
         .D(key_mem_new[31]), .Z(key_mem_0__127__N_6368[31])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i32_3_lut_4_lut.init = 16'hf2d0;
    PFUMX keylen_I_0_Mux_64_i1 (.BLUT(key_mem_new_127__N_7264[64]), .ALUT(prev_key1_new_127__N_7520[64]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[64])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    PFUMX i25891 (.BLUT(n8_adj_8868), .ALUT(n9_adj_8867), .C0(\muxed_round_nr[1] ), 
          .Z(n31050));
    LUT4 mux_12_i33_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [32]), 
         .D(key_mem_new[32]), .Z(key_mem_0__127__N_6368[32])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i33_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i34_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [33]), 
         .D(key_mem_new[33]), .Z(key_mem_0__127__N_6368[33])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i34_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i35_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [34]), 
         .D(key_mem_new[34]), .Z(key_mem_0__127__N_6368[34])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i35_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i36_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [35]), 
         .D(key_mem_new[35]), .Z(key_mem_0__127__N_6368[35])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i36_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i37_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [36]), 
         .D(key_mem_new[36]), .Z(key_mem_0__127__N_6368[36])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i37_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25221 (.BLUT(n8_adj_8866), .ALUT(n9_adj_8864), .C0(\muxed_round_nr[1] ), 
          .Z(n30380));
    LUT4 mux_12_i38_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [37]), 
         .D(key_mem_new[37]), .Z(key_mem_0__127__N_6368[37])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i38_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i39_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [38]), 
         .D(key_mem_new[38]), .Z(key_mem_0__127__N_6368[38])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i39_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i66_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [65]), 
         .D(key_mem_new[65]), .Z(key_mem_0__127__N_6368[65])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i66_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25896 (.BLUT(n1_adj_8863), .ALUT(n2_adj_8861), .C0(\muxed_round_nr[1] ), 
          .Z(n31055));
    PFUMX i25897 (.BLUT(n4_adj_8860), .ALUT(n5_adj_8859), .C0(\muxed_round_nr[1] ), 
          .Z(n31056));
    LUT4 mux_12_i67_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [66]), 
         .D(key_mem_new[66]), .Z(key_mem_0__127__N_6368[66])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i67_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25226 (.BLUT(n1_adj_8858), .ALUT(n2_adj_8856), .C0(\muxed_round_nr[1] ), 
          .Z(n30385));
    PFUMX i25898 (.BLUT(n8_adj_8857), .ALUT(n9_adj_8855), .C0(\muxed_round_nr[1] ), 
          .Z(n31057));
    LUT4 mux_12_i68_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [67]), 
         .D(key_mem_new[67]), .Z(key_mem_0__127__N_6368[67])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i68_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25227 (.BLUT(n4_adj_8853), .ALUT(n5_adj_8852), .C0(\muxed_round_nr[1] ), 
          .Z(n30386));
    LUT4 mux_12_i69_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [68]), 
         .D(key_mem_new[68]), .Z(key_mem_0__127__N_6368[68])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i69_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i70_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [69]), 
         .D(key_mem_new[69]), .Z(key_mem_0__127__N_6368[69])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i70_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25903 (.BLUT(n1_adj_8851), .ALUT(n2_adj_8850), .C0(\muxed_round_nr[1] ), 
          .Z(n31062));
    LUT4 mux_12_i71_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [70]), 
         .D(key_mem_new[70]), .Z(key_mem_0__127__N_6368[70])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i71_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25228 (.BLUT(n8_adj_8849), .ALUT(n9_adj_8846), .C0(\muxed_round_nr[1] ), 
          .Z(n30387));
    PFUMX i25904 (.BLUT(n4_adj_8848), .ALUT(n5_adj_8847), .C0(\muxed_round_nr[1] ), 
          .Z(n31063));
    LUT4 mux_12_i72_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [71]), 
         .D(key_mem_new[71]), .Z(key_mem_0__127__N_6368[71])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i72_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i73_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [72]), 
         .D(key_mem_new[72]), .Z(key_mem_0__127__N_6368[72])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i73_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i74_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [73]), 
         .D(key_mem_new[73]), .Z(key_mem_0__127__N_6368[73])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i74_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i75_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [74]), 
         .D(key_mem_new[74]), .Z(key_mem_0__127__N_6368[74])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i75_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25905 (.BLUT(n8_adj_8845), .ALUT(n9_adj_8843), .C0(\muxed_round_nr[1] ), 
          .Z(n31064));
    LUT4 mux_12_i76_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [75]), 
         .D(key_mem_new[75]), .Z(key_mem_0__127__N_6368[75])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i76_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i77_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [76]), 
         .D(key_mem_new[76]), .Z(key_mem_0__127__N_6368[76])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i77_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i78_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [77]), 
         .D(key_mem_new[77]), .Z(key_mem_0__127__N_6368[77])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i78_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25233 (.BLUT(n1_adj_8841), .ALUT(n2_adj_8839), .C0(\muxed_round_nr[1] ), 
          .Z(n30392));
    LUT4 mux_12_i79_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [78]), 
         .D(key_mem_new[78]), .Z(key_mem_0__127__N_6368[78])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i79_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25910 (.BLUT(n1_adj_8840), .ALUT(n2_adj_8838), .C0(\muxed_round_nr[1] ), 
          .Z(n31069));
    LUT4 mux_12_i80_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [79]), 
         .D(key_mem_new[79]), .Z(key_mem_0__127__N_6368[79])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i80_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25234 (.BLUT(n4_adj_8836), .ALUT(n5_adj_8834), .C0(\muxed_round_nr[1] ), 
          .Z(n30393));
    PFUMX i25911 (.BLUT(n4_adj_8837), .ALUT(n5_adj_8835), .C0(\muxed_round_nr[1] ), 
          .Z(n31070));
    PFUMX i25912 (.BLUT(n8_adj_8833), .ALUT(n9_adj_8832), .C0(\muxed_round_nr[1] ), 
          .Z(n31071));
    LUT4 mux_12_i81_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [80]), 
         .D(key_mem_new[80]), .Z(key_mem_0__127__N_6368[80])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i81_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25235 (.BLUT(n8_adj_8831), .ALUT(n9_adj_8830), .C0(\muxed_round_nr[1] ), 
          .Z(n30394));
    LUT4 mux_12_i82_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [81]), 
         .D(key_mem_new[81]), .Z(key_mem_0__127__N_6368[81])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i82_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i83_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [82]), 
         .D(key_mem_new[82]), .Z(key_mem_0__127__N_6368[82])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i83_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i84_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [83]), 
         .D(key_mem_new[83]), .Z(key_mem_0__127__N_6368[83])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i84_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i85_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [84]), 
         .D(key_mem_new[84]), .Z(key_mem_0__127__N_6368[84])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i85_3_lut_4_lut.init = 16'hf2d0;
    PFUMX keylen_I_0_Mux_119_i1 (.BLUT(key_mem_new_127__N_7264[119]), .ALUT(prev_key1_new_127__N_7520[119]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[119])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    LUT4 mux_12_i86_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [85]), 
         .D(key_mem_new[85]), .Z(key_mem_0__127__N_6368[85])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i86_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25240 (.BLUT(n1_adj_8827), .ALUT(n2_adj_8826), .C0(\muxed_round_nr[1] ), 
          .Z(n30399));
    LUT4 mux_12_i87_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [86]), 
         .D(key_mem_new[86]), .Z(key_mem_0__127__N_6368[86])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i87_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i88_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [87]), 
         .D(key_mem_new[87]), .Z(key_mem_0__127__N_6368[87])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i88_3_lut_4_lut.init = 16'hf2d0;
    PFUMX keylen_I_0_Mux_118_i1 (.BLUT(key_mem_new_127__N_7264[118]), .ALUT(prev_key1_new_127__N_7520[118]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[118])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    LUT4 mux_12_i89_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [88]), 
         .D(key_mem_new[88]), .Z(key_mem_0__127__N_6368[88])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i89_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i90_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [89]), 
         .D(key_mem_new[89]), .Z(key_mem_0__127__N_6368[89])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i90_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25917 (.BLUT(n1_adj_8824), .ALUT(n2_adj_8822), .C0(\muxed_round_nr[1] ), 
          .Z(n31076));
    PFUMX i25241 (.BLUT(n4_adj_8825), .ALUT(n5_adj_8823), .C0(\muxed_round_nr[1] ), 
          .Z(n30400));
    PFUMX keylen_I_0_Mux_117_i1 (.BLUT(key_mem_new_127__N_7264[117]), .ALUT(prev_key1_new_127__N_7520[117]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[117])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    LUT4 mux_12_i91_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [90]), 
         .D(key_mem_new[90]), .Z(key_mem_0__127__N_6368[90])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i91_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i92_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [91]), 
         .D(key_mem_new[91]), .Z(key_mem_0__127__N_6368[91])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i92_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25918 (.BLUT(n4_adj_8821), .ALUT(n5_adj_8818), .C0(\muxed_round_nr[1] ), 
          .Z(n31077));
    PFUMX keylen_I_0_Mux_116_i1 (.BLUT(key_mem_new_127__N_7264[116]), .ALUT(prev_key1_new_127__N_7520[116]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[116])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    LUT4 mux_12_i93_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [92]), 
         .D(key_mem_new[92]), .Z(key_mem_0__127__N_6368[92])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i93_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25242 (.BLUT(n8_adj_8820), .ALUT(n9_adj_8819), .C0(\muxed_round_nr[1] ), 
          .Z(n30401));
    LUT4 mux_12_i94_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [93]), 
         .D(key_mem_new[93]), .Z(key_mem_0__127__N_6368[93])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i94_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i95_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [94]), 
         .D(key_mem_new[94]), .Z(key_mem_0__127__N_6368[94])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i95_3_lut_4_lut.init = 16'hf2d0;
    PFUMX keylen_I_0_Mux_115_i1 (.BLUT(key_mem_new_127__N_7264[115]), .ALUT(prev_key1_new_127__N_7520[115]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[115])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    LUT4 mux_12_i96_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [95]), 
         .D(key_mem_new[95]), .Z(key_mem_0__127__N_6368[95])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i96_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i97_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [96]), 
         .D(key_mem_new[96]), .Z(key_mem_0__127__N_6368[96])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i97_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i98_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [97]), 
         .D(key_mem_new[97]), .Z(key_mem_0__127__N_6368[97])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i98_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25919 (.BLUT(n8_adj_8816), .ALUT(n9_adj_8814), .C0(\muxed_round_nr[1] ), 
          .Z(n31078));
    PFUMX i25247 (.BLUT(n1_adj_8815), .ALUT(n2_adj_8813), .C0(\muxed_round_nr[1] ), 
          .Z(n30406));
    PFUMX keylen_I_0_Mux_114_i1 (.BLUT(key_mem_new_127__N_7264[114]), .ALUT(prev_key1_new_127__N_7520[114]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[114])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    LUT4 mux_12_i99_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [98]), 
         .D(key_mem_new[98]), .Z(key_mem_0__127__N_6368[98])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i99_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i100_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [99]), 
         .D(key_mem_new[99]), .Z(key_mem_0__127__N_6368[99])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i100_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i101_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [100]), 
         .D(key_mem_new[100]), .Z(key_mem_0__127__N_6368[100])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i101_3_lut_4_lut.init = 16'hf2d0;
    PFUMX keylen_I_0_Mux_113_i1 (.BLUT(key_mem_new_127__N_7264[113]), .ALUT(prev_key1_new_127__N_7520[113]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[113])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    LUT4 mux_12_i102_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [101]), 
         .D(key_mem_new[101]), .Z(key_mem_0__127__N_6368[101])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i102_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i103_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [102]), 
         .D(key_mem_new[102]), .Z(key_mem_0__127__N_6368[102])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i103_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25248 (.BLUT(n4_adj_8812), .ALUT(n5_adj_8811), .C0(\muxed_round_nr[1] ), 
          .Z(n30407));
    PFUMX i25249 (.BLUT(n8_adj_8809), .ALUT(n9_adj_8808), .C0(\muxed_round_nr[1] ), 
          .Z(n30408));
    LUT4 mux_12_i104_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [103]), 
         .D(key_mem_new[103]), .Z(key_mem_0__127__N_6368[103])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i104_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i105_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [104]), 
         .D(key_mem_new[104]), .Z(key_mem_0__127__N_6368[104])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i105_3_lut_4_lut.init = 16'hf2d0;
    PFUMX keylen_I_0_Mux_112_i1 (.BLUT(key_mem_new_127__N_7264[112]), .ALUT(prev_key1_new_127__N_7520[112]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[112])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    LUT4 mux_12_i106_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [105]), 
         .D(key_mem_new[105]), .Z(key_mem_0__127__N_6368[105])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i106_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25254 (.BLUT(n1_adj_8806), .ALUT(n2_adj_8804), .C0(\muxed_round_nr[1] ), 
          .Z(n30413));
    LUT4 mux_12_i107_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [106]), 
         .D(key_mem_new[106]), .Z(key_mem_0__127__N_6368[106])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i107_3_lut_4_lut.init = 16'hf2d0;
    PFUMX keylen_I_0_Mux_111_i1 (.BLUT(key_mem_new_127__N_7264[111]), .ALUT(prev_key1_new_127__N_7520[111]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[111])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    PFUMX i25924 (.BLUT(n1_adj_8805), .ALUT(n2_adj_8803), .C0(\muxed_round_nr[1] ), 
          .Z(n31083));
    LUT4 mux_12_i108_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [107]), 
         .D(key_mem_new[107]), .Z(key_mem_0__127__N_6368[107])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i108_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i109_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [108]), 
         .D(key_mem_new[108]), .Z(key_mem_0__127__N_6368[108])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i109_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i110_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [109]), 
         .D(key_mem_new[109]), .Z(key_mem_0__127__N_6368[109])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i110_3_lut_4_lut.init = 16'hf2d0;
    PFUMX keylen_I_0_Mux_110_i1 (.BLUT(key_mem_new_127__N_7264[110]), .ALUT(prev_key1_new_127__N_7520[110]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[110])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    PFUMX i25255 (.BLUT(n4_adj_8801), .ALUT(n5_adj_8800), .C0(\muxed_round_nr[1] ), 
          .Z(n30414));
    PFUMX i25925 (.BLUT(n4_adj_8802), .ALUT(n5_adj_8798), .C0(\muxed_round_nr[1] ), 
          .Z(n31084));
    LUT4 mux_12_i111_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [110]), 
         .D(key_mem_new[110]), .Z(key_mem_0__127__N_6368[110])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i111_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i112_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [111]), 
         .D(key_mem_new[111]), .Z(key_mem_0__127__N_6368[111])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i112_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25256 (.BLUT(n8_adj_8799), .ALUT(n9_adj_8797), .C0(\muxed_round_nr[1] ), 
          .Z(n30415));
    PFUMX keylen_I_0_Mux_109_i1 (.BLUT(key_mem_new_127__N_7264[109]), .ALUT(prev_key1_new_127__N_7520[109]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[109])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    LUT4 mux_12_i113_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [112]), 
         .D(key_mem_new[112]), .Z(key_mem_0__127__N_6368[112])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i113_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i114_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [113]), 
         .D(key_mem_new[113]), .Z(key_mem_0__127__N_6368[113])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i114_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i115_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [114]), 
         .D(key_mem_new[114]), .Z(key_mem_0__127__N_6368[114])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i115_3_lut_4_lut.init = 16'hf2d0;
    PFUMX keylen_I_0_Mux_108_i1 (.BLUT(key_mem_new_127__N_7264[108]), .ALUT(prev_key1_new_127__N_7520[108]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[108])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    LUT4 mux_12_i116_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [115]), 
         .D(key_mem_new[115]), .Z(key_mem_0__127__N_6368[115])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i116_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i117_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [116]), 
         .D(key_mem_new[116]), .Z(key_mem_0__127__N_6368[116])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i117_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i118_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [117]), 
         .D(key_mem_new[117]), .Z(key_mem_0__127__N_6368[117])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i118_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25926 (.BLUT(n8_adj_8795), .ALUT(n9_adj_8794), .C0(\muxed_round_nr[1] ), 
          .Z(n31085));
    LUT4 mux_12_i119_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [118]), 
         .D(key_mem_new[118]), .Z(key_mem_0__127__N_6368[118])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i119_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i120_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [119]), 
         .D(key_mem_new[119]), .Z(key_mem_0__127__N_6368[119])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i120_3_lut_4_lut.init = 16'hf2d0;
    PFUMX keylen_I_0_Mux_107_i1 (.BLUT(key_mem_new_127__N_7264[107]), .ALUT(prev_key1_new_127__N_7520[107]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[107])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    PFUMX i25261 (.BLUT(n1_adj_8793), .ALUT(n2_adj_8792), .C0(\muxed_round_nr[1] ), 
          .Z(n30420));
    LUT4 mux_12_i121_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [120]), 
         .D(key_mem_new[120]), .Z(key_mem_0__127__N_6368[120])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i121_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i122_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [121]), 
         .D(key_mem_new[121]), .Z(key_mem_0__127__N_6368[121])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i122_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25262 (.BLUT(n4_adj_8791), .ALUT(n5_adj_8789), .C0(\muxed_round_nr[1] ), 
          .Z(n30421));
    PFUMX keylen_I_0_Mux_106_i1 (.BLUT(key_mem_new_127__N_7264[106]), .ALUT(prev_key1_new_127__N_7520[106]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[106])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    PFUMX i25263 (.BLUT(n8_adj_8788), .ALUT(n9_adj_8787), .C0(\muxed_round_nr[1] ), 
          .Z(n30422));
    LUT4 mux_12_i123_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [122]), 
         .D(key_mem_new[122]), .Z(key_mem_0__127__N_6368[122])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i123_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i124_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [123]), 
         .D(key_mem_new[123]), .Z(key_mem_0__127__N_6368[123])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i124_3_lut_4_lut.init = 16'hf2d0;
    PFUMX keylen_I_0_Mux_105_i1 (.BLUT(key_mem_new_127__N_7264[105]), .ALUT(prev_key1_new_127__N_7520[105]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[105])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    LUT4 mux_12_i125_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [124]), 
         .D(key_mem_new[124]), .Z(key_mem_0__127__N_6368[124])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i125_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25931 (.BLUT(n1_adj_8786), .ALUT(n2_adj_8785), .C0(\muxed_round_nr[1] ), 
          .Z(n31090));
    LUT4 mux_12_i126_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [125]), 
         .D(key_mem_new[125]), .Z(key_mem_0__127__N_6368[125])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i126_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i127_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [126]), 
         .D(key_mem_new[126]), .Z(key_mem_0__127__N_6368[126])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i127_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_12_i128_3_lut_4_lut (.A(n33938), .B(n33937), .C(\key_mem[11] [127]), 
         .D(key_mem_new[127]), .Z(key_mem_0__127__N_6368[127])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_12_i128_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_11_i65_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [64]), 
         .D(key_mem_new[64]), .Z(key_mem_0__127__N_6496[64])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i65_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i39_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [38]), 
         .D(key_mem_new[38]), .Z(key_mem_0__127__N_6496[38])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i39_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25932 (.BLUT(n4_adj_8783), .ALUT(n5_adj_8782), .C0(\muxed_round_nr[1] ), 
          .Z(n31091));
    PFUMX keylen_I_0_Mux_104_i1 (.BLUT(key_mem_new_127__N_7264[104]), .ALUT(prev_key1_new_127__N_7520[104]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[104])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    LUT4 mux_11_i40_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [39]), 
         .D(key_mem_new[39]), .Z(key_mem_0__127__N_6496[39])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i40_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i41_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [40]), 
         .D(key_mem_new[40]), .Z(key_mem_0__127__N_6496[40])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i41_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i42_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [41]), 
         .D(key_mem_new[41]), .Z(key_mem_0__127__N_6496[41])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i42_3_lut_4_lut.init = 16'hf4b0;
    PFUMX keylen_I_0_Mux_103_i1 (.BLUT(key_mem_new_127__N_7264[103]), .ALUT(prev_key1_new_127__N_7520[103]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[103])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    LUT4 mux_11_i43_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [42]), 
         .D(key_mem_new[42]), .Z(key_mem_0__127__N_6496[42])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i43_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25933 (.BLUT(n8_adj_8781), .ALUT(n9_adj_8780), .C0(\muxed_round_nr[1] ), 
          .Z(n31092));
    LUT4 mux_11_i44_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [43]), 
         .D(key_mem_new[43]), .Z(key_mem_0__127__N_6496[43])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i44_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25268 (.BLUT(n1_adj_8779), .ALUT(n2_adj_8778), .C0(\muxed_round_nr[1] ), 
          .Z(n30427));
    LUT4 mux_11_i45_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [44]), 
         .D(key_mem_new[44]), .Z(key_mem_0__127__N_6496[44])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i45_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i46_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [45]), 
         .D(key_mem_new[45]), .Z(key_mem_0__127__N_6496[45])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i46_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i47_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [46]), 
         .D(key_mem_new[46]), .Z(key_mem_0__127__N_6496[46])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i47_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25269 (.BLUT(n4_adj_8777), .ALUT(n5_adj_8776), .C0(\muxed_round_nr[1] ), 
          .Z(n30428));
    LUT4 mux_11_i48_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [47]), 
         .D(key_mem_new[47]), .Z(key_mem_0__127__N_6496[47])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i48_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i49_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [48]), 
         .D(key_mem_new[48]), .Z(key_mem_0__127__N_6496[48])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i49_3_lut_4_lut.init = 16'hf4b0;
    PFUMX keylen_I_0_Mux_102_i1 (.BLUT(key_mem_new_127__N_7264[102]), .ALUT(prev_key1_new_127__N_7520[102]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[102])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    LUT4 mux_11_i50_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [49]), 
         .D(key_mem_new[49]), .Z(key_mem_0__127__N_6496[49])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i50_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i51_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [50]), 
         .D(key_mem_new[50]), .Z(key_mem_0__127__N_6496[50])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i51_3_lut_4_lut.init = 16'hf4b0;
    PFUMX keylen_I_0_Mux_101_i1 (.BLUT(key_mem_new_127__N_7264[101]), .ALUT(prev_key1_new_127__N_7520[101]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[101])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    PFUMX i25270 (.BLUT(n8_adj_8774), .ALUT(n9_adj_8773), .C0(\muxed_round_nr[1] ), 
          .Z(n30429));
    LUT4 mux_11_i52_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [51]), 
         .D(key_mem_new[51]), .Z(key_mem_0__127__N_6496[51])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i52_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i53_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [52]), 
         .D(key_mem_new[52]), .Z(key_mem_0__127__N_6496[52])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i53_3_lut_4_lut.init = 16'hf4b0;
    PFUMX keylen_I_0_Mux_100_i1 (.BLUT(key_mem_new_127__N_7264[100]), .ALUT(prev_key1_new_127__N_7520[100]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[100])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    LUT4 mux_11_i54_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [53]), 
         .D(key_mem_new[53]), .Z(key_mem_0__127__N_6496[53])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i54_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i55_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [54]), 
         .D(key_mem_new[54]), .Z(key_mem_0__127__N_6496[54])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i55_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25938 (.BLUT(n1_adj_8772), .ALUT(n2_adj_8771), .C0(\muxed_round_nr[1] ), 
          .Z(n31097));
    PFUMX keylen_I_0_Mux_99_i1 (.BLUT(key_mem_new_127__N_7264[99]), .ALUT(prev_key1_new_127__N_7520[99]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[99])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    LUT4 mux_11_i56_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [55]), 
         .D(key_mem_new[55]), .Z(key_mem_0__127__N_6496[55])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i56_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i57_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [56]), 
         .D(key_mem_new[56]), .Z(key_mem_0__127__N_6496[56])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i57_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i58_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [57]), 
         .D(key_mem_new[57]), .Z(key_mem_0__127__N_6496[57])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i58_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i59_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [58]), 
         .D(key_mem_new[58]), .Z(key_mem_0__127__N_6496[58])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i59_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i60_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [59]), 
         .D(key_mem_new[59]), .Z(key_mem_0__127__N_6496[59])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i60_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i61_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [60]), 
         .D(key_mem_new[60]), .Z(key_mem_0__127__N_6496[60])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i61_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25939 (.BLUT(n4_adj_8769), .ALUT(n5_adj_8767), .C0(\muxed_round_nr[1] ), 
          .Z(n31098));
    PFUMX keylen_I_0_Mux_98_i1 (.BLUT(key_mem_new_127__N_7264[98]), .ALUT(prev_key1_new_127__N_7520[98]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[98])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    LUT4 mux_11_i62_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [61]), 
         .D(key_mem_new[61]), .Z(key_mem_0__127__N_6496[61])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i62_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i63_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [62]), 
         .D(key_mem_new[62]), .Z(key_mem_0__127__N_6496[62])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i63_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i64_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [63]), 
         .D(key_mem_new[63]), .Z(key_mem_0__127__N_6496[63])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i64_3_lut_4_lut.init = 16'hf4b0;
    PFUMX keylen_I_0_Mux_97_i1 (.BLUT(key_mem_new_127__N_7264[97]), .ALUT(prev_key1_new_127__N_7520[97]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[97])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    LUT4 mux_11_i1_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [0]), 
         .D(key_mem_new[0]), .Z(key_mem_0__127__N_6496[0])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i1_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25275 (.BLUT(n1_adj_8768), .ALUT(n2_adj_8766), .C0(\muxed_round_nr[1] ), 
          .Z(n30434));
    PFUMX i25940 (.BLUT(n8_adj_8765), .ALUT(n9_adj_8762), .C0(\muxed_round_nr[1] ), 
          .Z(n31099));
    LUT4 mux_11_i2_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [1]), 
         .D(key_mem_new[1]), .Z(key_mem_0__127__N_6496[1])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i2_3_lut_4_lut.init = 16'hf4b0;
    PFUMX keylen_I_0_Mux_96_i1 (.BLUT(key_mem_new_127__N_7264[96]), .ALUT(prev_key1_new_127__N_7520[96]), 
          .C0(\key_mem_ctrl.num_rounds[2] ), .Z(prev_key1_new_127__N_4787[96])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=15, LSE_RCOL=22, LSE_LLINE=151, LSE_RLINE=165 */ ;
    LUT4 mux_11_i3_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [2]), 
         .D(key_mem_new[2]), .Z(key_mem_0__127__N_6496[2])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i3_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i4_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [3]), 
         .D(key_mem_new[3]), .Z(key_mem_0__127__N_6496[3])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i4_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25276 (.BLUT(n4_adj_8764), .ALUT(n5_adj_8763), .C0(\muxed_round_nr[1] ), 
          .Z(n30435));
    LUT4 mux_11_i5_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [4]), 
         .D(key_mem_new[4]), .Z(key_mem_0__127__N_6496[4])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i5_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25277 (.BLUT(n8_adj_8760), .ALUT(n9_adj_8759), .C0(\muxed_round_nr[1] ), 
          .Z(n30436));
    LUT4 mux_11_i6_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [5]), 
         .D(key_mem_new[5]), .Z(key_mem_0__127__N_6496[5])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i6_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i7_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [6]), 
         .D(key_mem_new[6]), .Z(key_mem_0__127__N_6496[6])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i7_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i8_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [7]), 
         .D(key_mem_new[7]), .Z(key_mem_0__127__N_6496[7])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i8_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i9_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [8]), 
         .D(key_mem_new[8]), .Z(key_mem_0__127__N_6496[8])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i9_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i10_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [9]), 
         .D(key_mem_new[9]), .Z(key_mem_0__127__N_6496[9])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i10_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25945 (.BLUT(n1_adj_8757), .ALUT(n2_adj_8755), .C0(\muxed_round_nr[1] ), 
          .Z(n31104));
    LUT4 mux_11_i11_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [10]), 
         .D(key_mem_new[10]), .Z(key_mem_0__127__N_6496[10])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i11_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25282 (.BLUT(n1_adj_8756), .ALUT(n2_adj_8754), .C0(\muxed_round_nr[1] ), 
          .Z(n30441));
    LUT4 mux_11_i12_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [11]), 
         .D(key_mem_new[11]), .Z(key_mem_0__127__N_6496[11])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i12_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25946 (.BLUT(n4_adj_8753), .ALUT(n5_adj_8752), .C0(\muxed_round_nr[1] ), 
          .Z(n31105));
    LUT4 mux_11_i13_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [12]), 
         .D(key_mem_new[12]), .Z(key_mem_0__127__N_6496[12])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i13_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25283 (.BLUT(n4_adj_8751), .ALUT(n5_adj_8748), .C0(\muxed_round_nr[1] ), 
          .Z(n30442));
    LUT4 mux_11_i14_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [13]), 
         .D(key_mem_new[13]), .Z(key_mem_0__127__N_6496[13])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i14_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25947 (.BLUT(n8_adj_8750), .ALUT(n9_adj_8749), .C0(\muxed_round_nr[1] ), 
          .Z(n31106));
    LUT4 mux_11_i15_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [14]), 
         .D(key_mem_new[14]), .Z(key_mem_0__127__N_6496[14])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i15_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i16_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [15]), 
         .D(key_mem_new[15]), .Z(key_mem_0__127__N_6496[15])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i16_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25284 (.BLUT(n8_adj_8747), .ALUT(n9_adj_8746), .C0(\muxed_round_nr[1] ), 
          .Z(n30443));
    LUT4 mux_11_i17_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [16]), 
         .D(key_mem_new[16]), .Z(key_mem_0__127__N_6496[16])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i17_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i18_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [17]), 
         .D(key_mem_new[17]), .Z(key_mem_0__127__N_6496[17])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i18_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i19_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [18]), 
         .D(key_mem_new[18]), .Z(key_mem_0__127__N_6496[18])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i19_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i20_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [19]), 
         .D(key_mem_new[19]), .Z(key_mem_0__127__N_6496[19])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i20_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25289 (.BLUT(n1_adj_8743), .ALUT(n2_adj_8742), .C0(\muxed_round_nr[1] ), 
          .Z(n30448));
    LUT4 mux_11_i21_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [20]), 
         .D(key_mem_new[20]), .Z(key_mem_0__127__N_6496[20])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i21_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i22_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [21]), 
         .D(key_mem_new[21]), .Z(key_mem_0__127__N_6496[21])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i22_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25952 (.BLUT(n1_adj_8741), .ALUT(n2_adj_8740), .C0(\muxed_round_nr[1] ), 
          .Z(n31111));
    LUT4 mux_11_i23_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [22]), 
         .D(key_mem_new[22]), .Z(key_mem_0__127__N_6496[22])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i23_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25953 (.BLUT(n4_adj_8739), .ALUT(n5_adj_8737), .C0(\muxed_round_nr[1] ), 
          .Z(n31112));
    PFUMX i25290 (.BLUT(n4_adj_8738), .ALUT(n5_adj_8736), .C0(\muxed_round_nr[1] ), 
          .Z(n30449));
    LUT4 mux_11_i24_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [23]), 
         .D(key_mem_new[23]), .Z(key_mem_0__127__N_6496[23])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i24_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25954 (.BLUT(n8_adj_8735), .ALUT(n9_adj_8733), .C0(\muxed_round_nr[1] ), 
          .Z(n31113));
    PFUMX i25291 (.BLUT(n8_adj_8734), .ALUT(n9_adj_8732), .C0(\muxed_round_nr[1] ), 
          .Z(n30450));
    LUT4 mux_11_i25_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [24]), 
         .D(key_mem_new[24]), .Z(key_mem_0__127__N_6496[24])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i25_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i26_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [25]), 
         .D(key_mem_new[25]), .Z(key_mem_0__127__N_6496[25])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i26_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i27_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [26]), 
         .D(key_mem_new[26]), .Z(key_mem_0__127__N_6496[26])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i27_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i28_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [27]), 
         .D(key_mem_new[27]), .Z(key_mem_0__127__N_6496[27])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i28_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i29_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [28]), 
         .D(key_mem_new[28]), .Z(key_mem_0__127__N_6496[28])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i29_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25296 (.BLUT(n1_adj_8729), .ALUT(n2_adj_8727), .C0(\muxed_round_nr[1] ), 
          .Z(n30455));
    PFUMX i25959 (.BLUT(n1_adj_8728), .ALUT(n2_adj_8726), .C0(\muxed_round_nr[1] ), 
          .Z(n31118));
    LUT4 mux_11_i30_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [29]), 
         .D(key_mem_new[29]), .Z(key_mem_0__127__N_6496[29])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i30_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25297 (.BLUT(n4_adj_8725), .ALUT(n5_adj_8724), .C0(\muxed_round_nr[1] ), 
          .Z(n30456));
    LUT4 mux_11_i31_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [30]), 
         .D(key_mem_new[30]), .Z(key_mem_0__127__N_6496[30])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i31_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25298 (.BLUT(n8_adj_8723), .ALUT(n9_adj_8722), .C0(\muxed_round_nr[1] ), 
          .Z(n30457));
    PFUMX i25960 (.BLUT(n4_adj_8720), .ALUT(n5_adj_8719), .C0(\muxed_round_nr[1] ), 
          .Z(n31119));
    LUT4 mux_11_i32_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [31]), 
         .D(key_mem_new[31]), .Z(key_mem_0__127__N_6496[31])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i32_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25961 (.BLUT(n8_adj_8718), .ALUT(n9_adj_8717), .C0(\muxed_round_nr[1] ), 
          .Z(n31120));
    LUT4 mux_11_i33_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [32]), 
         .D(key_mem_new[32]), .Z(key_mem_0__127__N_6496[32])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i33_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25303 (.BLUT(n1_adj_8715), .ALUT(n2_adj_8714), .C0(\muxed_round_nr[1] ), 
          .Z(n30462));
    LUT4 mux_11_i34_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [33]), 
         .D(key_mem_new[33]), .Z(key_mem_0__127__N_6496[33])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i34_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i35_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [34]), 
         .D(key_mem_new[34]), .Z(key_mem_0__127__N_6496[34])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i35_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25966 (.BLUT(n1_adj_8712), .ALUT(n2_adj_8706), .C0(\muxed_round_nr[1] ), 
          .Z(n31125));
    LUT4 mux_11_i36_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [35]), 
         .D(key_mem_new[35]), .Z(key_mem_0__127__N_6496[35])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i36_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25304 (.BLUT(n4_adj_8713), .ALUT(n5_adj_8711), .C0(\muxed_round_nr[1] ), 
          .Z(n30463));
    LUT4 mux_11_i37_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [36]), 
         .D(key_mem_new[36]), .Z(key_mem_0__127__N_6496[36])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i37_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25305 (.BLUT(n8_adj_8710), .ALUT(n9_adj_8707), .C0(\muxed_round_nr[1] ), 
          .Z(n30464));
    LUT4 mux_11_i38_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [37]), 
         .D(key_mem_new[37]), .Z(key_mem_0__127__N_6496[37])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i38_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i66_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [65]), 
         .D(key_mem_new[65]), .Z(key_mem_0__127__N_6496[65])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i66_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i67_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [66]), 
         .D(key_mem_new[66]), .Z(key_mem_0__127__N_6496[66])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i67_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25967 (.BLUT(n4_adj_8705), .ALUT(n5_adj_8703), .C0(\muxed_round_nr[1] ), 
          .Z(n31126));
    LUT4 mux_11_i68_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [67]), 
         .D(key_mem_new[67]), .Z(key_mem_0__127__N_6496[67])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i68_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25310 (.BLUT(n1_adj_8683), .ALUT(n2_adj_8680), .C0(\muxed_round_nr[1] ), 
          .Z(n30469));
    PFUMX i25968 (.BLUT(n8_adj_8682), .ALUT(n9_adj_8681), .C0(\muxed_round_nr[1] ), 
          .Z(n31127));
    LUT4 mux_11_i69_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [68]), 
         .D(key_mem_new[68]), .Z(key_mem_0__127__N_6496[68])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i69_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25311 (.BLUT(n4_adj_8678), .ALUT(n5_adj_8677), .C0(\muxed_round_nr[1] ), 
          .Z(n30470));
    LUT4 mux_11_i70_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [69]), 
         .D(key_mem_new[69]), .Z(key_mem_0__127__N_6496[69])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i70_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i71_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [70]), 
         .D(key_mem_new[70]), .Z(key_mem_0__127__N_6496[70])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i71_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i72_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [71]), 
         .D(key_mem_new[71]), .Z(key_mem_0__127__N_6496[71])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i72_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25973 (.BLUT(n1_adj_8674), .ALUT(n2_adj_8670), .C0(\muxed_round_nr[1] ), 
          .Z(n31132));
    LUT4 mux_11_i73_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [72]), 
         .D(key_mem_new[72]), .Z(key_mem_0__127__N_6496[72])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i73_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25312 (.BLUT(n8_adj_8673), .ALUT(n9_adj_8672), .C0(\muxed_round_nr[1] ), 
          .Z(n30471));
    LUT4 mux_11_i74_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [73]), 
         .D(key_mem_new[73]), .Z(key_mem_0__127__N_6496[73])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i74_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i75_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [74]), 
         .D(key_mem_new[74]), .Z(key_mem_0__127__N_6496[74])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i75_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25974 (.BLUT(n4_adj_8668), .ALUT(n5_adj_8666), .C0(\muxed_round_nr[1] ), 
          .Z(n31133));
    LUT4 mux_11_i76_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [75]), 
         .D(key_mem_new[75]), .Z(key_mem_0__127__N_6496[75])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i76_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25317 (.BLUT(n1_adj_8669), .ALUT(n2_adj_8667), .C0(\muxed_round_nr[1] ), 
          .Z(n30476));
    LUT4 mux_11_i77_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [76]), 
         .D(key_mem_new[76]), .Z(key_mem_0__127__N_6496[76])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i77_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25318 (.BLUT(n4_adj_8665), .ALUT(n5_adj_8664), .C0(\muxed_round_nr[1] ), 
          .Z(n30477));
    PFUMX i25975 (.BLUT(n8_adj_8663), .ALUT(n9_adj_8661), .C0(\muxed_round_nr[1] ), 
          .Z(n31134));
    PFUMX i25319 (.BLUT(n8_adj_8662), .ALUT(n9_adj_8660), .C0(\muxed_round_nr[1] ), 
          .Z(n30478));
    LUT4 mux_11_i78_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [77]), 
         .D(key_mem_new[77]), .Z(key_mem_0__127__N_6496[77])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i78_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i79_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [78]), 
         .D(key_mem_new[78]), .Z(key_mem_0__127__N_6496[78])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i79_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i80_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [79]), 
         .D(key_mem_new[79]), .Z(key_mem_0__127__N_6496[79])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i80_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i81_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [80]), 
         .D(key_mem_new[80]), .Z(key_mem_0__127__N_6496[80])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i81_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i82_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [81]), 
         .D(key_mem_new[81]), .Z(key_mem_0__127__N_6496[81])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i82_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i83_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [82]), 
         .D(key_mem_new[82]), .Z(key_mem_0__127__N_6496[82])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i83_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25324 (.BLUT(n1_adj_8657), .ALUT(n2_adj_8656), .C0(\muxed_round_nr[1] ), 
          .Z(n30483));
    LUT4 mux_11_i84_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [83]), 
         .D(key_mem_new[83]), .Z(key_mem_0__127__N_6496[83])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i84_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i85_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [84]), 
         .D(key_mem_new[84]), .Z(key_mem_0__127__N_6496[84])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i85_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25325 (.BLUT(n4_adj_8655), .ALUT(n5_adj_8654), .C0(\muxed_round_nr[1] ), 
          .Z(n30484));
    LUT4 mux_11_i86_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [85]), 
         .D(key_mem_new[85]), .Z(key_mem_0__127__N_6496[85])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i86_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i87_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [86]), 
         .D(key_mem_new[86]), .Z(key_mem_0__127__N_6496[86])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i87_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25326 (.BLUT(n8_adj_8653), .ALUT(n9_adj_8652), .C0(\muxed_round_nr[1] ), 
          .Z(n30485));
    LUT4 mux_11_i88_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [87]), 
         .D(key_mem_new[87]), .Z(key_mem_0__127__N_6496[87])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i88_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i89_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [88]), 
         .D(key_mem_new[88]), .Z(key_mem_0__127__N_6496[88])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i89_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i90_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [89]), 
         .D(key_mem_new[89]), .Z(key_mem_0__127__N_6496[89])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i90_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i91_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [90]), 
         .D(key_mem_new[90]), .Z(key_mem_0__127__N_6496[90])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i91_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i92_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [91]), 
         .D(key_mem_new[91]), .Z(key_mem_0__127__N_6496[91])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i92_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i93_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [92]), 
         .D(key_mem_new[92]), .Z(key_mem_0__127__N_6496[92])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i93_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25331 (.BLUT(n1_adj_8643), .ALUT(n2_adj_8638), .C0(\muxed_round_nr[1] ), 
          .Z(n30490));
    LUT4 mux_11_i94_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [93]), 
         .D(key_mem_new[93]), .Z(key_mem_0__127__N_6496[93])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i94_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i95_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [94]), 
         .D(key_mem_new[94]), .Z(key_mem_0__127__N_6496[94])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i95_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25332 (.BLUT(n4_adj_8635), .ALUT(n5_adj_8634), .C0(\muxed_round_nr[1] ), 
          .Z(n30491));
    LUT4 mux_11_i96_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [95]), 
         .D(key_mem_new[95]), .Z(key_mem_0__127__N_6496[95])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i96_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i97_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [96]), 
         .D(key_mem_new[96]), .Z(key_mem_0__127__N_6496[96])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i97_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25333 (.BLUT(n8_adj_8632), .ALUT(n9_adj_8631), .C0(\muxed_round_nr[1] ), 
          .Z(n30492));
    LUT4 mux_11_i98_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [97]), 
         .D(key_mem_new[97]), .Z(key_mem_0__127__N_6496[97])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i98_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i99_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [98]), 
         .D(key_mem_new[98]), .Z(key_mem_0__127__N_6496[98])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i99_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i100_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [99]), 
         .D(key_mem_new[99]), .Z(key_mem_0__127__N_6496[99])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i100_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i101_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [100]), 
         .D(key_mem_new[100]), .Z(key_mem_0__127__N_6496[100])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i101_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i102_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [101]), 
         .D(key_mem_new[101]), .Z(key_mem_0__127__N_6496[101])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i102_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i103_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [102]), 
         .D(key_mem_new[102]), .Z(key_mem_0__127__N_6496[102])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i103_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25338 (.BLUT(n1_adj_8629), .ALUT(n2_adj_8628), .C0(\muxed_round_nr[1] ), 
          .Z(n30497));
    LUT4 mux_11_i104_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [103]), 
         .D(key_mem_new[103]), .Z(key_mem_0__127__N_6496[103])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i104_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i105_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [104]), 
         .D(key_mem_new[104]), .Z(key_mem_0__127__N_6496[104])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i105_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i106_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [105]), 
         .D(key_mem_new[105]), .Z(key_mem_0__127__N_6496[105])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i106_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25339 (.BLUT(n4_adj_8624), .ALUT(n5_adj_8623), .C0(\muxed_round_nr[1] ), 
          .Z(n30498));
    LUT4 mux_11_i107_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [106]), 
         .D(key_mem_new[106]), .Z(key_mem_0__127__N_6496[106])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i107_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i108_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [107]), 
         .D(key_mem_new[107]), .Z(key_mem_0__127__N_6496[107])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i108_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25340 (.BLUT(n8_adj_8621), .ALUT(n9_adj_8619), .C0(\muxed_round_nr[1] ), 
          .Z(n30499));
    LUT4 mux_11_i109_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [108]), 
         .D(key_mem_new[108]), .Z(key_mem_0__127__N_6496[108])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i109_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i110_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [109]), 
         .D(key_mem_new[109]), .Z(key_mem_0__127__N_6496[109])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i110_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i111_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [110]), 
         .D(key_mem_new[110]), .Z(key_mem_0__127__N_6496[110])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i111_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i112_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [111]), 
         .D(key_mem_new[111]), .Z(key_mem_0__127__N_6496[111])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i112_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25345 (.BLUT(n1_adj_8613), .ALUT(n2_adj_8612), .C0(\muxed_round_nr[1] ), 
          .Z(n30504));
    LUT4 mux_11_i113_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [112]), 
         .D(key_mem_new[112]), .Z(key_mem_0__127__N_6496[112])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i113_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25346 (.BLUT(n4_adj_8610), .ALUT(n5_adj_8609), .C0(\muxed_round_nr[1] ), 
          .Z(n30505));
    LUT4 mux_11_i114_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [113]), 
         .D(key_mem_new[113]), .Z(key_mem_0__127__N_6496[113])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i114_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i115_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [114]), 
         .D(key_mem_new[114]), .Z(key_mem_0__127__N_6496[114])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i115_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i116_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [115]), 
         .D(key_mem_new[115]), .Z(key_mem_0__127__N_6496[115])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i116_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25347 (.BLUT(n8_adj_8606), .ALUT(n9_adj_8605), .C0(\muxed_round_nr[1] ), 
          .Z(n30506));
    LUT4 mux_11_i117_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [116]), 
         .D(key_mem_new[116]), .Z(key_mem_0__127__N_6496[116])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i117_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i118_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [117]), 
         .D(key_mem_new[117]), .Z(key_mem_0__127__N_6496[117])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i118_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i119_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [118]), 
         .D(key_mem_new[118]), .Z(key_mem_0__127__N_6496[118])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i119_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i120_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [119]), 
         .D(key_mem_new[119]), .Z(key_mem_0__127__N_6496[119])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i120_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25352 (.BLUT(n1_adj_8597), .ALUT(n2_adj_8595), .C0(\muxed_round_nr[1] ), 
          .Z(n30511));
    LUT4 mux_11_i121_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [120]), 
         .D(key_mem_new[120]), .Z(key_mem_0__127__N_6496[120])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i121_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25353 (.BLUT(n4_adj_8594), .ALUT(n5_adj_8593), .C0(\muxed_round_nr[1] ), 
          .Z(n30512));
    LUT4 mux_11_i122_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [121]), 
         .D(key_mem_new[121]), .Z(key_mem_0__127__N_6496[121])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i122_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25354 (.BLUT(n8_adj_8592), .ALUT(n9_adj_8591), .C0(\muxed_round_nr[1] ), 
          .Z(n30513));
    LUT4 mux_11_i123_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [122]), 
         .D(key_mem_new[122]), .Z(key_mem_0__127__N_6496[122])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i123_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i124_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [123]), 
         .D(key_mem_new[123]), .Z(key_mem_0__127__N_6496[123])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i124_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i125_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [124]), 
         .D(key_mem_new[124]), .Z(key_mem_0__127__N_6496[124])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i125_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i126_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [125]), 
         .D(key_mem_new[125]), .Z(key_mem_0__127__N_6496[125])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i126_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i127_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [126]), 
         .D(key_mem_new[126]), .Z(key_mem_0__127__N_6496[126])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i127_3_lut_4_lut.init = 16'hf4b0;
    FD1P3AX key_mem_ctrl_reg_FSM_i0_i2 (.D(n33951), .SP(key_mem_ctrl_we), 
            .CK(clk_c), .Q(n6361[2]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam key_mem_ctrl_reg_FSM_i0_i2.GSR = "ENABLED";
    FD1P3AY key_mem_ctrl_reg_FSM_i0_i3 (.D(n28834), .SP(key_mem_ctrl_we), 
            .CK(clk_c), .Q(n6361[3]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam key_mem_ctrl_reg_FSM_i0_i3.GSR = "ENABLED";
    LUT4 mux_11_i128_3_lut_4_lut (.A(n33943), .B(n33911), .C(\key_mem[12] [127]), 
         .D(key_mem_new[127]), .Z(key_mem_0__127__N_6496[127])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_11_i128_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25359 (.BLUT(n1_adj_8585), .ALUT(n2_adj_8584), .C0(\muxed_round_nr[1] ), 
          .Z(n30518));
    PFUMX i25360 (.BLUT(n4_adj_8583), .ALUT(n5_adj_8582), .C0(\muxed_round_nr[1] ), 
          .Z(n30519));
    LUT4 mux_10_i65_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [64]), 
         .D(key_mem_new[64]), .Z(key_mem_0__127__N_6624[64])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i65_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i39_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [38]), 
         .D(key_mem_new[38]), .Z(key_mem_0__127__N_6624[38])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i39_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i40_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [39]), 
         .D(key_mem_new[39]), .Z(key_mem_0__127__N_6624[39])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i40_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i41_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [40]), 
         .D(key_mem_new[40]), .Z(key_mem_0__127__N_6624[40])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i41_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25361 (.BLUT(n8_adj_8580), .ALUT(n9_adj_8579), .C0(\muxed_round_nr[1] ), 
          .Z(n30520));
    LUT4 mux_10_i42_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [41]), 
         .D(key_mem_new[41]), .Z(key_mem_0__127__N_6624[41])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i42_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i43_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [42]), 
         .D(key_mem_new[42]), .Z(key_mem_0__127__N_6624[42])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i43_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i44_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [43]), 
         .D(key_mem_new[43]), .Z(key_mem_0__127__N_6624[43])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i44_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i45_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [44]), 
         .D(key_mem_new[44]), .Z(key_mem_0__127__N_6624[44])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i45_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i46_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [45]), 
         .D(key_mem_new[45]), .Z(key_mem_0__127__N_6624[45])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i46_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i47_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [46]), 
         .D(key_mem_new[46]), .Z(key_mem_0__127__N_6624[46])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i47_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i48_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [47]), 
         .D(key_mem_new[47]), .Z(key_mem_0__127__N_6624[47])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i48_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i49_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [48]), 
         .D(key_mem_new[48]), .Z(key_mem_0__127__N_6624[48])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i49_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i50_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [49]), 
         .D(key_mem_new[49]), .Z(key_mem_0__127__N_6624[49])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i50_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i51_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [50]), 
         .D(key_mem_new[50]), .Z(key_mem_0__127__N_6624[50])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i51_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i52_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [51]), 
         .D(key_mem_new[51]), .Z(key_mem_0__127__N_6624[51])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i52_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i53_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [52]), 
         .D(key_mem_new[52]), .Z(key_mem_0__127__N_6624[52])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i53_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i54_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [53]), 
         .D(key_mem_new[53]), .Z(key_mem_0__127__N_6624[53])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i54_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i55_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [54]), 
         .D(key_mem_new[54]), .Z(key_mem_0__127__N_6624[54])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i55_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i56_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [55]), 
         .D(key_mem_new[55]), .Z(key_mem_0__127__N_6624[55])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i56_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i57_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [56]), 
         .D(key_mem_new[56]), .Z(key_mem_0__127__N_6624[56])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i57_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i58_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [57]), 
         .D(key_mem_new[57]), .Z(key_mem_0__127__N_6624[57])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i58_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i59_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [58]), 
         .D(key_mem_new[58]), .Z(key_mem_0__127__N_6624[58])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i59_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i60_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [59]), 
         .D(key_mem_new[59]), .Z(key_mem_0__127__N_6624[59])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i60_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i61_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [60]), 
         .D(key_mem_new[60]), .Z(key_mem_0__127__N_6624[60])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i61_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i62_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [61]), 
         .D(key_mem_new[61]), .Z(key_mem_0__127__N_6624[61])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i62_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i63_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [62]), 
         .D(key_mem_new[62]), .Z(key_mem_0__127__N_6624[62])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i63_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25366 (.BLUT(n1_adj_8576), .ALUT(n2_adj_8575), .C0(\muxed_round_nr[1] ), 
          .Z(n30525));
    LUT4 mux_10_i64_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [63]), 
         .D(key_mem_new[63]), .Z(key_mem_0__127__N_6624[63])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i64_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i1_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [0]), 
         .D(key_mem_new[0]), .Z(key_mem_0__127__N_6624[0])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i1_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i2_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [1]), 
         .D(key_mem_new[1]), .Z(key_mem_0__127__N_6624[1])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i2_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i3_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [2]), 
         .D(key_mem_new[2]), .Z(key_mem_0__127__N_6624[2])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i3_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i4_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [3]), 
         .D(key_mem_new[3]), .Z(key_mem_0__127__N_6624[3])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i4_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i5_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [4]), 
         .D(key_mem_new[4]), .Z(key_mem_0__127__N_6624[4])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i5_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i6_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [5]), 
         .D(key_mem_new[5]), .Z(key_mem_0__127__N_6624[5])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i6_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i7_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [6]), 
         .D(key_mem_new[6]), .Z(key_mem_0__127__N_6624[6])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i7_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i8_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [7]), 
         .D(key_mem_new[7]), .Z(key_mem_0__127__N_6624[7])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i8_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i9_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [8]), 
         .D(key_mem_new[8]), .Z(key_mem_0__127__N_6624[8])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i9_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i10_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [9]), 
         .D(key_mem_new[9]), .Z(key_mem_0__127__N_6624[9])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i10_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i11_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [10]), 
         .D(key_mem_new[10]), .Z(key_mem_0__127__N_6624[10])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i11_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i12_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [11]), 
         .D(key_mem_new[11]), .Z(key_mem_0__127__N_6624[11])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i12_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25367 (.BLUT(n4_adj_8574), .ALUT(n5_adj_8573), .C0(\muxed_round_nr[1] ), 
          .Z(n30526));
    LUT4 mux_10_i13_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [12]), 
         .D(key_mem_new[12]), .Z(key_mem_0__127__N_6624[12])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i13_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i14_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [13]), 
         .D(key_mem_new[13]), .Z(key_mem_0__127__N_6624[13])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i14_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i15_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [14]), 
         .D(key_mem_new[14]), .Z(key_mem_0__127__N_6624[14])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i15_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i16_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [15]), 
         .D(key_mem_new[15]), .Z(key_mem_0__127__N_6624[15])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i16_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i17_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [16]), 
         .D(key_mem_new[16]), .Z(key_mem_0__127__N_6624[16])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i17_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i18_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [17]), 
         .D(key_mem_new[17]), .Z(key_mem_0__127__N_6624[17])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i18_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25368 (.BLUT(n8_adj_8572), .ALUT(n9_adj_8571), .C0(\muxed_round_nr[1] ), 
          .Z(n30527));
    LUT4 mux_10_i19_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [18]), 
         .D(key_mem_new[18]), .Z(key_mem_0__127__N_6624[18])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i19_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i20_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [19]), 
         .D(key_mem_new[19]), .Z(key_mem_0__127__N_6624[19])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i20_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i21_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [20]), 
         .D(key_mem_new[20]), .Z(key_mem_0__127__N_6624[20])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i21_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i22_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [21]), 
         .D(key_mem_new[21]), .Z(key_mem_0__127__N_6624[21])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i22_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i23_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [22]), 
         .D(key_mem_new[22]), .Z(key_mem_0__127__N_6624[22])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i23_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i24_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [23]), 
         .D(key_mem_new[23]), .Z(key_mem_0__127__N_6624[23])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i24_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i25_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [24]), 
         .D(key_mem_new[24]), .Z(key_mem_0__127__N_6624[24])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i25_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i26_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [25]), 
         .D(key_mem_new[25]), .Z(key_mem_0__127__N_6624[25])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i26_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i27_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [26]), 
         .D(key_mem_new[26]), .Z(key_mem_0__127__N_6624[26])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i27_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i28_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [27]), 
         .D(key_mem_new[27]), .Z(key_mem_0__127__N_6624[27])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i28_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i29_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [28]), 
         .D(key_mem_new[28]), .Z(key_mem_0__127__N_6624[28])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i29_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i30_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [29]), 
         .D(key_mem_new[29]), .Z(key_mem_0__127__N_6624[29])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i30_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i31_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [30]), 
         .D(key_mem_new[30]), .Z(key_mem_0__127__N_6624[30])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i31_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i32_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [31]), 
         .D(key_mem_new[31]), .Z(key_mem_0__127__N_6624[31])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i32_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i33_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [32]), 
         .D(key_mem_new[32]), .Z(key_mem_0__127__N_6624[32])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i33_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i34_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [33]), 
         .D(key_mem_new[33]), .Z(key_mem_0__127__N_6624[33])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i34_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i35_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [34]), 
         .D(key_mem_new[34]), .Z(key_mem_0__127__N_6624[34])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i35_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i36_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [35]), 
         .D(key_mem_new[35]), .Z(key_mem_0__127__N_6624[35])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i36_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i37_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [36]), 
         .D(key_mem_new[36]), .Z(key_mem_0__127__N_6624[36])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i37_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i38_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [37]), 
         .D(key_mem_new[37]), .Z(key_mem_0__127__N_6624[37])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i38_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i66_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [65]), 
         .D(key_mem_new[65]), .Z(key_mem_0__127__N_6624[65])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i66_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i67_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [66]), 
         .D(key_mem_new[66]), .Z(key_mem_0__127__N_6624[66])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i67_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i68_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [67]), 
         .D(key_mem_new[67]), .Z(key_mem_0__127__N_6624[67])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i68_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i69_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [68]), 
         .D(key_mem_new[68]), .Z(key_mem_0__127__N_6624[68])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i69_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i70_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [69]), 
         .D(key_mem_new[69]), .Z(key_mem_0__127__N_6624[69])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i70_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i71_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [70]), 
         .D(key_mem_new[70]), .Z(key_mem_0__127__N_6624[70])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i71_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25373 (.BLUT(n1_adj_8566), .ALUT(n2_adj_8565), .C0(\muxed_round_nr[1] ), 
          .Z(n30532));
    LUT4 mux_10_i72_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [71]), 
         .D(key_mem_new[71]), .Z(key_mem_0__127__N_6624[71])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i72_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i73_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [72]), 
         .D(key_mem_new[72]), .Z(key_mem_0__127__N_6624[72])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i73_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i74_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [73]), 
         .D(key_mem_new[73]), .Z(key_mem_0__127__N_6624[73])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i74_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i75_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [74]), 
         .D(key_mem_new[74]), .Z(key_mem_0__127__N_6624[74])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i75_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i76_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [75]), 
         .D(key_mem_new[75]), .Z(key_mem_0__127__N_6624[75])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i76_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i77_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [76]), 
         .D(key_mem_new[76]), .Z(key_mem_0__127__N_6624[76])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i77_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i78_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [77]), 
         .D(key_mem_new[77]), .Z(key_mem_0__127__N_6624[77])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i78_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i79_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [78]), 
         .D(key_mem_new[78]), .Z(key_mem_0__127__N_6624[78])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i79_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25374 (.BLUT(n4_adj_8561), .ALUT(n5_adj_8559), .C0(\muxed_round_nr[1] ), 
          .Z(n30533));
    LUT4 mux_10_i80_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [79]), 
         .D(key_mem_new[79]), .Z(key_mem_0__127__N_6624[79])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i80_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i81_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [80]), 
         .D(key_mem_new[80]), .Z(key_mem_0__127__N_6624[80])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i81_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i82_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [81]), 
         .D(key_mem_new[81]), .Z(key_mem_0__127__N_6624[81])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i82_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i83_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [82]), 
         .D(key_mem_new[82]), .Z(key_mem_0__127__N_6624[82])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i83_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i84_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [83]), 
         .D(key_mem_new[83]), .Z(key_mem_0__127__N_6624[83])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i84_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i85_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [84]), 
         .D(key_mem_new[84]), .Z(key_mem_0__127__N_6624[84])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i85_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i86_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [85]), 
         .D(key_mem_new[85]), .Z(key_mem_0__127__N_6624[85])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i86_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i87_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [86]), 
         .D(key_mem_new[86]), .Z(key_mem_0__127__N_6624[86])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i87_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i88_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [87]), 
         .D(key_mem_new[87]), .Z(key_mem_0__127__N_6624[87])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i88_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i89_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [88]), 
         .D(key_mem_new[88]), .Z(key_mem_0__127__N_6624[88])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i89_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i90_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [89]), 
         .D(key_mem_new[89]), .Z(key_mem_0__127__N_6624[89])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i90_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25375 (.BLUT(n8_adj_8558), .ALUT(n9_adj_8557), .C0(\muxed_round_nr[1] ), 
          .Z(n30534));
    LUT4 mux_10_i91_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [90]), 
         .D(key_mem_new[90]), .Z(key_mem_0__127__N_6624[90])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i91_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i92_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [91]), 
         .D(key_mem_new[91]), .Z(key_mem_0__127__N_6624[91])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i92_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i93_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [92]), 
         .D(key_mem_new[92]), .Z(key_mem_0__127__N_6624[92])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i93_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i94_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [93]), 
         .D(key_mem_new[93]), .Z(key_mem_0__127__N_6624[93])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i94_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i95_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [94]), 
         .D(key_mem_new[94]), .Z(key_mem_0__127__N_6624[94])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i95_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i96_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [95]), 
         .D(key_mem_new[95]), .Z(key_mem_0__127__N_6624[95])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i96_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i97_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [96]), 
         .D(key_mem_new[96]), .Z(key_mem_0__127__N_6624[96])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i97_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i98_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [97]), 
         .D(key_mem_new[97]), .Z(key_mem_0__127__N_6624[97])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i98_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i99_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [98]), 
         .D(key_mem_new[98]), .Z(key_mem_0__127__N_6624[98])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i99_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i100_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [99]), 
         .D(key_mem_new[99]), .Z(key_mem_0__127__N_6624[99])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i100_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i101_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [100]), 
         .D(key_mem_new[100]), .Z(key_mem_0__127__N_6624[100])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i101_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i102_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [101]), 
         .D(key_mem_new[101]), .Z(key_mem_0__127__N_6624[101])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i102_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i103_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [102]), 
         .D(key_mem_new[102]), .Z(key_mem_0__127__N_6624[102])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i103_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i104_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [103]), 
         .D(key_mem_new[103]), .Z(key_mem_0__127__N_6624[103])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i104_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i105_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [104]), 
         .D(key_mem_new[104]), .Z(key_mem_0__127__N_6624[104])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i105_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i106_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [105]), 
         .D(key_mem_new[105]), .Z(key_mem_0__127__N_6624[105])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i106_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i107_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [106]), 
         .D(key_mem_new[106]), .Z(key_mem_0__127__N_6624[106])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i107_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i108_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [107]), 
         .D(key_mem_new[107]), .Z(key_mem_0__127__N_6624[107])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i108_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i109_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [108]), 
         .D(key_mem_new[108]), .Z(key_mem_0__127__N_6624[108])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i109_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25380 (.BLUT(n1_adj_8554), .ALUT(n2_adj_8553), .C0(\muxed_round_nr[1] ), 
          .Z(n30539));
    LUT4 mux_10_i110_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [109]), 
         .D(key_mem_new[109]), .Z(key_mem_0__127__N_6624[109])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i110_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i111_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [110]), 
         .D(key_mem_new[110]), .Z(key_mem_0__127__N_6624[110])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i111_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i112_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [111]), 
         .D(key_mem_new[111]), .Z(key_mem_0__127__N_6624[111])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i112_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i113_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [112]), 
         .D(key_mem_new[112]), .Z(key_mem_0__127__N_6624[112])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i113_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i114_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [113]), 
         .D(key_mem_new[113]), .Z(key_mem_0__127__N_6624[113])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i114_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i115_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [114]), 
         .D(key_mem_new[114]), .Z(key_mem_0__127__N_6624[114])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i115_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i116_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [115]), 
         .D(key_mem_new[115]), .Z(key_mem_0__127__N_6624[115])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i116_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i117_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [116]), 
         .D(key_mem_new[116]), .Z(key_mem_0__127__N_6624[116])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i117_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i118_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [117]), 
         .D(key_mem_new[117]), .Z(key_mem_0__127__N_6624[117])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i118_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i119_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [118]), 
         .D(key_mem_new[118]), .Z(key_mem_0__127__N_6624[118])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i119_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i120_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [119]), 
         .D(key_mem_new[119]), .Z(key_mem_0__127__N_6624[119])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i120_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i121_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [120]), 
         .D(key_mem_new[120]), .Z(key_mem_0__127__N_6624[120])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i121_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i122_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [121]), 
         .D(key_mem_new[121]), .Z(key_mem_0__127__N_6624[121])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i122_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i123_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [122]), 
         .D(key_mem_new[122]), .Z(key_mem_0__127__N_6624[122])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i123_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i124_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [123]), 
         .D(key_mem_new[123]), .Z(key_mem_0__127__N_6624[123])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i124_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i125_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [124]), 
         .D(key_mem_new[124]), .Z(key_mem_0__127__N_6624[124])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i125_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i25381 (.BLUT(n4_adj_8552), .ALUT(n5_adj_8551), .C0(\muxed_round_nr[1] ), 
          .Z(n30540));
    LUT4 mux_10_i126_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [125]), 
         .D(key_mem_new[125]), .Z(key_mem_0__127__N_6624[125])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i126_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i127_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [126]), 
         .D(key_mem_new[126]), .Z(key_mem_0__127__N_6624[126])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i127_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i128_3_lut_4_lut (.A(n33945), .B(n33911), .C(\key_mem[13] [127]), 
         .D(key_mem_new[127]), .Z(key_mem_0__127__N_6624[127])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam mux_10_i128_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_85_i120_3_lut_rep_287_4_lut (.A(n33945), .B(n33944), .C(n4_adj_8421), 
         .D(\key_reg[4] [23]), .Z(n33591)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_85_i120_3_lut_rep_287_4_lut.init = 16'hf1e0;
    PFUMX i25382 (.BLUT(n8_adj_8547), .ALUT(n9_adj_8546), .C0(\muxed_round_nr[1] ), 
          .Z(n30541));
    LUT4 mux_85_i97_3_lut_rep_310_4_lut (.A(n33945), .B(n33944), .C(n8487), 
         .D(\key_reg[4] [0]), .Z(n33614)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_85_i97_3_lut_rep_310_4_lut.init = 16'hf1e0;
    LUT4 mux_85_i98_3_lut_rep_309_4_lut (.A(n33945), .B(n33944), .C(n8929), 
         .D(\key_reg[4] [1]), .Z(n33613)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_85_i98_3_lut_rep_309_4_lut.init = 16'hf1e0;
    LUT4 mux_85_i99_3_lut_rep_308_4_lut (.A(n33945), .B(n33944), .C(n4_adj_8332), 
         .D(\key_reg[4] [2]), .Z(n33612)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_85_i99_3_lut_rep_308_4_lut.init = 16'hf1e0;
    LUT4 mux_85_i100_3_lut_rep_307_4_lut (.A(n33945), .B(n33944), .C(n4_adj_8333), 
         .D(\key_reg[4] [3]), .Z(n33611)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_85_i100_3_lut_rep_307_4_lut.init = 16'hf1e0;
    LUT4 mux_85_i101_3_lut_rep_306_4_lut (.A(n33945), .B(n33944), .C(n4_adj_8335), 
         .D(\key_reg[4] [4]), .Z(n33610)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_85_i101_3_lut_rep_306_4_lut.init = 16'hf1e0;
    LUT4 mux_85_i102_3_lut_rep_305_4_lut (.A(n33945), .B(n33944), .C(n4_adj_8336), 
         .D(\key_reg[4] [5]), .Z(n33609)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_85_i102_3_lut_rep_305_4_lut.init = 16'hf1e0;
    LUT4 mux_85_i103_3_lut_rep_304_4_lut (.A(n33945), .B(n33944), .C(n4_adj_8337), 
         .D(\key_reg[4] [6]), .Z(n33608)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_85_i103_3_lut_rep_304_4_lut.init = 16'hf1e0;
    LUT4 mux_85_i104_3_lut_rep_303_4_lut (.A(n33945), .B(n33944), .C(n4_adj_8339), 
         .D(\key_reg[4] [7]), .Z(n33607)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_85_i104_3_lut_rep_303_4_lut.init = 16'hf1e0;
    LUT4 mux_85_i105_3_lut_rep_302_4_lut (.A(n33945), .B(n33944), .C(n4_adj_8343), 
         .D(\key_reg[4] [8]), .Z(n33606)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_85_i105_3_lut_rep_302_4_lut.init = 16'hf1e0;
    LUT4 mux_85_i106_3_lut_rep_301_4_lut (.A(n33945), .B(n33944), .C(n4_adj_8349), 
         .D(\key_reg[4] [9]), .Z(n33605)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_85_i106_3_lut_rep_301_4_lut.init = 16'hf1e0;
    LUT4 mux_85_i107_3_lut_rep_300_4_lut (.A(n33945), .B(n33944), .C(n4), 
         .D(\key_reg[4] [10]), .Z(n33604)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_85_i107_3_lut_rep_300_4_lut.init = 16'hf1e0;
    LUT4 mux_85_i108_3_lut_rep_299_4_lut (.A(n33945), .B(n33944), .C(n4_adj_8361), 
         .D(\key_reg[4] [11]), .Z(n33603)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_85_i108_3_lut_rep_299_4_lut.init = 16'hf1e0;
    LUT4 mux_85_i109_3_lut_rep_298_4_lut (.A(n33945), .B(n33944), .C(n4_adj_8367), 
         .D(\key_reg[4] [12]), .Z(n33602)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_85_i109_3_lut_rep_298_4_lut.init = 16'hf1e0;
    LUT4 mux_85_i110_3_lut_rep_297_4_lut (.A(n33945), .B(n33944), .C(n4_adj_8373), 
         .D(\key_reg[4] [13]), .Z(n33601)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_85_i110_3_lut_rep_297_4_lut.init = 16'hf1e0;
    LUT4 mux_85_i111_3_lut_rep_296_4_lut (.A(n33945), .B(n33944), .C(n4_adj_8377), 
         .D(\key_reg[4] [14]), .Z(n33600)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_85_i111_3_lut_rep_296_4_lut.init = 16'hf1e0;
    LUT4 mux_85_i112_3_lut_rep_295_4_lut (.A(n33945), .B(n33944), .C(n4_adj_8381), 
         .D(\key_reg[4] [15]), .Z(n33599)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_85_i112_3_lut_rep_295_4_lut.init = 16'hf1e0;
    LUT4 mux_85_i113_3_lut_rep_294_4_lut (.A(n33945), .B(n33944), .C(n4_adj_8386), 
         .D(\key_reg[4] [16]), .Z(n33598)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_85_i113_3_lut_rep_294_4_lut.init = 16'hf1e0;
    LUT4 mux_85_i114_3_lut_rep_293_4_lut (.A(n33945), .B(n33944), .C(n4_adj_8390), 
         .D(\key_reg[4] [17]), .Z(n33597)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_85_i114_3_lut_rep_293_4_lut.init = 16'hf1e0;
    LUT4 mux_85_i115_3_lut_rep_292_4_lut (.A(n33945), .B(n33944), .C(n4_adj_8395), 
         .D(\key_reg[4] [18]), .Z(n33596)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_85_i115_3_lut_rep_292_4_lut.init = 16'hf1e0;
    LUT4 mux_85_i116_3_lut_rep_291_4_lut (.A(n33945), .B(n33944), .C(n4_adj_8400), 
         .D(\key_reg[4] [19]), .Z(n33595)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_85_i116_3_lut_rep_291_4_lut.init = 16'hf1e0;
    LUT4 mux_85_i117_3_lut_rep_290_4_lut (.A(n33945), .B(n33944), .C(n4_adj_8403), 
         .D(\key_reg[4] [20]), .Z(n33594)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_85_i117_3_lut_rep_290_4_lut.init = 16'hf1e0;
    LUT4 mux_85_i118_3_lut_rep_289_4_lut (.A(n33945), .B(n33944), .C(n4_adj_8410), 
         .D(\key_reg[4] [21]), .Z(n33593)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_85_i118_3_lut_rep_289_4_lut.init = 16'hf1e0;
    LUT4 mux_85_i119_3_lut_rep_288_4_lut (.A(n33945), .B(n33944), .C(n4_adj_8417), 
         .D(\key_reg[4] [22]), .Z(n33592)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_85_i119_3_lut_rep_288_4_lut.init = 16'hf1e0;
    LUT4 mux_85_i128_3_lut_rep_222_4_lut (.A(n33945), .B(n33944), .C(n4_adj_8457), 
         .D(\key_reg[4] [31]), .Z(n33526)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_85_i128_3_lut_rep_222_4_lut.init = 16'hf1e0;
    LUT4 mux_85_i127_3_lut_rep_223_4_lut (.A(n33945), .B(n33944), .C(n4_adj_8455), 
         .D(\key_reg[4] [30]), .Z(n33527)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_85_i127_3_lut_rep_223_4_lut.init = 16'hf1e0;
    LUT4 mux_85_i126_3_lut_rep_224_4_lut (.A(n33945), .B(n33944), .C(n4_adj_8451), 
         .D(\key_reg[4] [29]), .Z(n33528)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_85_i126_3_lut_rep_224_4_lut.init = 16'hf1e0;
    LUT4 mux_85_i125_3_lut_rep_225_4_lut (.A(n33945), .B(n33944), .C(n4_adj_8449), 
         .D(\key_reg[4] [28]), .Z(n33529)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_85_i125_3_lut_rep_225_4_lut.init = 16'hf1e0;
    LUT4 mux_85_i124_3_lut_rep_226_4_lut (.A(n33945), .B(n33944), .C(n4_adj_8444), 
         .D(\key_reg[4] [27]), .Z(n33530)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_85_i124_3_lut_rep_226_4_lut.init = 16'hf1e0;
    LUT4 mux_85_i123_3_lut_rep_227_4_lut (.A(n33945), .B(n33944), .C(n4_adj_8438), 
         .D(\key_reg[4] [26]), .Z(n33531)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_85_i123_3_lut_rep_227_4_lut.init = 16'hf1e0;
    LUT4 mux_85_i122_3_lut_rep_228_4_lut (.A(n33945), .B(n33944), .C(n4_adj_8430), 
         .D(\key_reg[4] [25]), .Z(n33532)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_85_i122_3_lut_rep_228_4_lut.init = 16'hf1e0;
    LUT4 mux_85_i121_3_lut_rep_229_4_lut (.A(n33945), .B(n33944), .C(n4_adj_8428), 
         .D(\key_reg[4] [24]), .Z(n33533)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_85_i121_3_lut_rep_229_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i1_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [0]), 
         .D(key_mem_new[0]), .Z(key_mem_0__127__N_5088[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i2_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [1]), 
         .D(key_mem_new[1]), .Z(key_mem_0__127__N_5088[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i3_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [2]), 
         .D(key_mem_new[2]), .Z(key_mem_0__127__N_5088[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i4_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [3]), 
         .D(key_mem_new[3]), .Z(key_mem_0__127__N_5088[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i5_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [4]), 
         .D(key_mem_new[4]), .Z(key_mem_0__127__N_5088[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i5_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25387 (.BLUT(n1_adj_8543), .ALUT(n2_adj_8541), .C0(\muxed_round_nr[1] ), 
          .Z(n30546));
    LUT4 mux_22_i6_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [5]), 
         .D(key_mem_new[5]), .Z(key_mem_0__127__N_5088[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i7_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [6]), 
         .D(key_mem_new[6]), .Z(key_mem_0__127__N_5088[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i8_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [7]), 
         .D(key_mem_new[7]), .Z(key_mem_0__127__N_5088[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i9_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [8]), 
         .D(key_mem_new[8]), .Z(key_mem_0__127__N_5088[8])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i9_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i10_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [9]), 
         .D(key_mem_new[9]), .Z(key_mem_0__127__N_5088[9])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i10_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i11_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [10]), 
         .D(key_mem_new[10]), .Z(key_mem_0__127__N_5088[10])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i11_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i12_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [11]), 
         .D(key_mem_new[11]), .Z(key_mem_0__127__N_5088[11])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i12_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i13_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [12]), 
         .D(key_mem_new[12]), .Z(key_mem_0__127__N_5088[12])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i13_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i14_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [13]), 
         .D(key_mem_new[13]), .Z(key_mem_0__127__N_5088[13])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i14_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i15_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [14]), 
         .D(key_mem_new[14]), .Z(key_mem_0__127__N_5088[14])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i15_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i16_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [15]), 
         .D(key_mem_new[15]), .Z(key_mem_0__127__N_5088[15])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i16_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i17_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [16]), 
         .D(key_mem_new[16]), .Z(key_mem_0__127__N_5088[16])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i17_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i18_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [17]), 
         .D(key_mem_new[17]), .Z(key_mem_0__127__N_5088[17])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i18_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i19_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [18]), 
         .D(key_mem_new[18]), .Z(key_mem_0__127__N_5088[18])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i19_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i20_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [19]), 
         .D(key_mem_new[19]), .Z(key_mem_0__127__N_5088[19])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i20_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i21_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [20]), 
         .D(key_mem_new[20]), .Z(key_mem_0__127__N_5088[20])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i21_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i22_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [21]), 
         .D(key_mem_new[21]), .Z(key_mem_0__127__N_5088[21])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i22_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i23_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [22]), 
         .D(key_mem_new[22]), .Z(key_mem_0__127__N_5088[22])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i23_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i24_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [23]), 
         .D(key_mem_new[23]), .Z(key_mem_0__127__N_5088[23])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i24_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i25_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [24]), 
         .D(key_mem_new[24]), .Z(key_mem_0__127__N_5088[24])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i25_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25388 (.BLUT(n4_adj_8540), .ALUT(n5_adj_8539), .C0(\muxed_round_nr[1] ), 
          .Z(n30547));
    LUT4 mux_22_i26_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [25]), 
         .D(key_mem_new[25]), .Z(key_mem_0__127__N_5088[25])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i26_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i27_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [26]), 
         .D(key_mem_new[26]), .Z(key_mem_0__127__N_5088[26])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i27_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i28_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [27]), 
         .D(key_mem_new[27]), .Z(key_mem_0__127__N_5088[27])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i28_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i29_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [28]), 
         .D(key_mem_new[28]), .Z(key_mem_0__127__N_5088[28])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i29_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i30_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [29]), 
         .D(key_mem_new[29]), .Z(key_mem_0__127__N_5088[29])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i30_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i31_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [30]), 
         .D(key_mem_new[30]), .Z(key_mem_0__127__N_5088[30])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i31_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i32_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [31]), 
         .D(key_mem_new[31]), .Z(key_mem_0__127__N_5088[31])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i32_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i33_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [32]), 
         .D(key_mem_new[32]), .Z(key_mem_0__127__N_5088[32])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i33_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i34_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [33]), 
         .D(key_mem_new[33]), .Z(key_mem_0__127__N_5088[33])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i34_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i35_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [34]), 
         .D(key_mem_new[34]), .Z(key_mem_0__127__N_5088[34])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i35_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i36_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [35]), 
         .D(key_mem_new[35]), .Z(key_mem_0__127__N_5088[35])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i36_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i37_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [36]), 
         .D(key_mem_new[36]), .Z(key_mem_0__127__N_5088[36])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i37_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i38_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [37]), 
         .D(key_mem_new[37]), .Z(key_mem_0__127__N_5088[37])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i38_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i39_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [38]), 
         .D(key_mem_new[38]), .Z(key_mem_0__127__N_5088[38])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i39_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i40_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [39]), 
         .D(key_mem_new[39]), .Z(key_mem_0__127__N_5088[39])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i40_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i41_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [40]), 
         .D(key_mem_new[40]), .Z(key_mem_0__127__N_5088[40])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i41_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25389 (.BLUT(n8_adj_8538), .ALUT(n9_adj_8537), .C0(\muxed_round_nr[1] ), 
          .Z(n30548));
    LUT4 mux_22_i42_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [41]), 
         .D(key_mem_new[41]), .Z(key_mem_0__127__N_5088[41])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i42_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i43_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [42]), 
         .D(key_mem_new[42]), .Z(key_mem_0__127__N_5088[42])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i43_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i44_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [43]), 
         .D(key_mem_new[43]), .Z(key_mem_0__127__N_5088[43])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i44_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i45_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [44]), 
         .D(key_mem_new[44]), .Z(key_mem_0__127__N_5088[44])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i45_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i46_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [45]), 
         .D(key_mem_new[45]), .Z(key_mem_0__127__N_5088[45])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i46_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i47_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [46]), 
         .D(key_mem_new[46]), .Z(key_mem_0__127__N_5088[46])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i47_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i48_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [47]), 
         .D(key_mem_new[47]), .Z(key_mem_0__127__N_5088[47])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i48_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i49_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [48]), 
         .D(key_mem_new[48]), .Z(key_mem_0__127__N_5088[48])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i49_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i50_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [49]), 
         .D(key_mem_new[49]), .Z(key_mem_0__127__N_5088[49])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i50_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i51_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [50]), 
         .D(key_mem_new[50]), .Z(key_mem_0__127__N_5088[50])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i51_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i52_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [51]), 
         .D(key_mem_new[51]), .Z(key_mem_0__127__N_5088[51])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i52_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i53_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [52]), 
         .D(key_mem_new[52]), .Z(key_mem_0__127__N_5088[52])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i53_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i54_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [53]), 
         .D(key_mem_new[53]), .Z(key_mem_0__127__N_5088[53])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i54_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i55_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [54]), 
         .D(key_mem_new[54]), .Z(key_mem_0__127__N_5088[54])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i55_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i56_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [55]), 
         .D(key_mem_new[55]), .Z(key_mem_0__127__N_5088[55])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i56_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i57_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [56]), 
         .D(key_mem_new[56]), .Z(key_mem_0__127__N_5088[56])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i57_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i58_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [57]), 
         .D(key_mem_new[57]), .Z(key_mem_0__127__N_5088[57])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i58_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i59_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [58]), 
         .D(key_mem_new[58]), .Z(key_mem_0__127__N_5088[58])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i59_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i60_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [59]), 
         .D(key_mem_new[59]), .Z(key_mem_0__127__N_5088[59])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i60_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i61_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [60]), 
         .D(key_mem_new[60]), .Z(key_mem_0__127__N_5088[60])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i61_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i62_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [61]), 
         .D(key_mem_new[61]), .Z(key_mem_0__127__N_5088[61])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i62_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i63_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [62]), 
         .D(key_mem_new[62]), .Z(key_mem_0__127__N_5088[62])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i63_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i64_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [63]), 
         .D(key_mem_new[63]), .Z(key_mem_0__127__N_5088[63])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i64_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i65_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [64]), 
         .D(key_mem_new[64]), .Z(key_mem_0__127__N_5088[64])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i65_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i66_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [65]), 
         .D(key_mem_new[65]), .Z(key_mem_0__127__N_5088[65])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i66_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i67_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [66]), 
         .D(key_mem_new[66]), .Z(key_mem_0__127__N_5088[66])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i67_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i68_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [67]), 
         .D(key_mem_new[67]), .Z(key_mem_0__127__N_5088[67])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i68_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i69_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [68]), 
         .D(key_mem_new[68]), .Z(key_mem_0__127__N_5088[68])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i69_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i70_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [69]), 
         .D(key_mem_new[69]), .Z(key_mem_0__127__N_5088[69])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i70_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i71_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [70]), 
         .D(key_mem_new[70]), .Z(key_mem_0__127__N_5088[70])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i71_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i72_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [71]), 
         .D(key_mem_new[71]), .Z(key_mem_0__127__N_5088[71])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i72_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i73_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [72]), 
         .D(key_mem_new[72]), .Z(key_mem_0__127__N_5088[72])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i73_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i74_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [73]), 
         .D(key_mem_new[73]), .Z(key_mem_0__127__N_5088[73])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i74_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i75_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [74]), 
         .D(key_mem_new[74]), .Z(key_mem_0__127__N_5088[74])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i75_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i76_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [75]), 
         .D(key_mem_new[75]), .Z(key_mem_0__127__N_5088[75])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i76_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i77_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [76]), 
         .D(key_mem_new[76]), .Z(key_mem_0__127__N_5088[76])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i77_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i78_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [77]), 
         .D(key_mem_new[77]), .Z(key_mem_0__127__N_5088[77])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i78_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i79_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [78]), 
         .D(key_mem_new[78]), .Z(key_mem_0__127__N_5088[78])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i79_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i80_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [79]), 
         .D(key_mem_new[79]), .Z(key_mem_0__127__N_5088[79])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i80_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i81_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [80]), 
         .D(key_mem_new[80]), .Z(key_mem_0__127__N_5088[80])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i81_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i82_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [81]), 
         .D(key_mem_new[81]), .Z(key_mem_0__127__N_5088[81])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i82_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i83_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [82]), 
         .D(key_mem_new[82]), .Z(key_mem_0__127__N_5088[82])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i83_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i84_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [83]), 
         .D(key_mem_new[83]), .Z(key_mem_0__127__N_5088[83])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i84_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i85_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [84]), 
         .D(key_mem_new[84]), .Z(key_mem_0__127__N_5088[84])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i85_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i86_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [85]), 
         .D(key_mem_new[85]), .Z(key_mem_0__127__N_5088[85])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i86_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i87_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [86]), 
         .D(key_mem_new[86]), .Z(key_mem_0__127__N_5088[86])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i87_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i88_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [87]), 
         .D(key_mem_new[87]), .Z(key_mem_0__127__N_5088[87])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i88_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i89_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [88]), 
         .D(key_mem_new[88]), .Z(key_mem_0__127__N_5088[88])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i89_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25394 (.BLUT(n1_adj_8533), .ALUT(n2_adj_8532), .C0(\muxed_round_nr[1] ), 
          .Z(n30553));
    LUT4 mux_22_i90_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [89]), 
         .D(key_mem_new[89]), .Z(key_mem_0__127__N_5088[89])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i90_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i91_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [90]), 
         .D(key_mem_new[90]), .Z(key_mem_0__127__N_5088[90])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i91_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i92_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [91]), 
         .D(key_mem_new[91]), .Z(key_mem_0__127__N_5088[91])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i92_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i93_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [92]), 
         .D(key_mem_new[92]), .Z(key_mem_0__127__N_5088[92])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i93_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i10 (.BLUT(n2531[0]), .ALUT(n8532), .C0(n29504), .Z(n10));
    LUT4 mux_22_i94_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [93]), 
         .D(key_mem_new[93]), .Z(key_mem_0__127__N_5088[93])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i94_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i95_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [94]), 
         .D(key_mem_new[94]), .Z(key_mem_0__127__N_5088[94])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i95_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i96_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [95]), 
         .D(key_mem_new[95]), .Z(key_mem_0__127__N_5088[95])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i96_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i97_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [96]), 
         .D(key_mem_new[96]), .Z(key_mem_0__127__N_5088[96])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i97_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i98_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [97]), 
         .D(key_mem_new[97]), .Z(key_mem_0__127__N_5088[97])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i98_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i99_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [98]), 
         .D(key_mem_new[98]), .Z(key_mem_0__127__N_5088[98])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i99_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i100_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [99]), 
         .D(key_mem_new[99]), .Z(key_mem_0__127__N_5088[99])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i100_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i101_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [100]), 
         .D(key_mem_new[100]), .Z(key_mem_0__127__N_5088[100])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i101_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i102_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [101]), 
         .D(key_mem_new[101]), .Z(key_mem_0__127__N_5088[101])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i102_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i103_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [102]), 
         .D(key_mem_new[102]), .Z(key_mem_0__127__N_5088[102])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i103_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i104_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [103]), 
         .D(key_mem_new[103]), .Z(key_mem_0__127__N_5088[103])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i104_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i105_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [104]), 
         .D(key_mem_new[104]), .Z(key_mem_0__127__N_5088[104])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i105_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i106_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [105]), 
         .D(key_mem_new[105]), .Z(key_mem_0__127__N_5088[105])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i106_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i107_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [106]), 
         .D(key_mem_new[106]), .Z(key_mem_0__127__N_5088[106])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i107_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i108_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [107]), 
         .D(key_mem_new[107]), .Z(key_mem_0__127__N_5088[107])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i108_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i109_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [108]), 
         .D(key_mem_new[108]), .Z(key_mem_0__127__N_5088[108])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i109_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i110_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [109]), 
         .D(key_mem_new[109]), .Z(key_mem_0__127__N_5088[109])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i110_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i111_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [110]), 
         .D(key_mem_new[110]), .Z(key_mem_0__127__N_5088[110])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i111_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i112_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [111]), 
         .D(key_mem_new[111]), .Z(key_mem_0__127__N_5088[111])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i112_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i113_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [112]), 
         .D(key_mem_new[112]), .Z(key_mem_0__127__N_5088[112])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i113_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i10_adj_664 (.BLUT(n2531[1]), .ALUT(n9616), .C0(n29504), .Z(n10_adj_8587));
    LUT4 mux_22_i114_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [113]), 
         .D(key_mem_new[113]), .Z(key_mem_0__127__N_5088[113])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i114_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i115_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [114]), 
         .D(key_mem_new[114]), .Z(key_mem_0__127__N_5088[114])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i115_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i116_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [115]), 
         .D(key_mem_new[115]), .Z(key_mem_0__127__N_5088[115])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i116_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i117_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [116]), 
         .D(key_mem_new[116]), .Z(key_mem_0__127__N_5088[116])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i117_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i118_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [117]), 
         .D(key_mem_new[117]), .Z(key_mem_0__127__N_5088[117])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i118_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i119_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [118]), 
         .D(key_mem_new[118]), .Z(key_mem_0__127__N_5088[118])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i119_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i120_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [119]), 
         .D(key_mem_new[119]), .Z(key_mem_0__127__N_5088[119])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i120_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i121_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [120]), 
         .D(key_mem_new[120]), .Z(key_mem_0__127__N_5088[120])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i121_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i122_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [121]), 
         .D(key_mem_new[121]), .Z(key_mem_0__127__N_5088[121])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i122_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i123_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [122]), 
         .D(key_mem_new[122]), .Z(key_mem_0__127__N_5088[122])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i123_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25395 (.BLUT(n4_adj_8531), .ALUT(n5_adj_8530), .C0(\muxed_round_nr[1] ), 
          .Z(n30554));
    LUT4 mux_22_i124_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [123]), 
         .D(key_mem_new[123]), .Z(key_mem_0__127__N_5088[123])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i124_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i125_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [124]), 
         .D(key_mem_new[124]), .Z(key_mem_0__127__N_5088[124])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i125_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i126_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [125]), 
         .D(key_mem_new[125]), .Z(key_mem_0__127__N_5088[125])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i126_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i127_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [126]), 
         .D(key_mem_new[126]), .Z(key_mem_0__127__N_5088[126])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i127_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i128_3_lut_4_lut (.A(n33945), .B(n33944), .C(\key_mem[1] [127]), 
         .D(key_mem_new[127]), .Z(key_mem_0__127__N_5088[127])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(264[26:44])
    defparam mux_22_i128_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i10_adj_665 (.BLUT(n2531[2]), .ALUT(n9618), .C0(n29504), .Z(n10_adj_8590));
    LUT4 mux_51_i81_3_lut_4_lut (.A(n33943), .B(n33944), .C(n33731), .D(\key_reg[1] [16]), 
         .Z(key_mem_new_127__N_7264[80])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_51_i81_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_51_i84_3_lut_4_lut (.A(n33943), .B(n33944), .C(n33728), .D(\key_reg[1] [19]), 
         .Z(key_mem_new_127__N_7264[83])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_51_i84_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_51_i85_3_lut_4_lut (.A(n33943), .B(n33944), .C(n33727), .D(\key_reg[1] [20]), 
         .Z(key_mem_new_127__N_7264[84])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_51_i85_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_51_i94_3_lut_4_lut (.A(n33943), .B(n33944), .C(n33615), .D(\key_reg[1] [29]), 
         .Z(key_mem_new_127__N_7264[93])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_51_i94_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_51_i93_3_lut_4_lut (.A(n33943), .B(n33944), .C(n33616), .D(\key_reg[1] [28]), 
         .Z(key_mem_new_127__N_7264[92])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_51_i93_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_51_i91_3_lut_4_lut (.A(n33943), .B(n33944), .C(n33618), .D(\key_reg[1] [26]), 
         .Z(key_mem_new_127__N_7264[90])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_51_i91_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_51_i89_3_lut_4_lut (.A(n33943), .B(n33944), .C(n33619), .D(\key_reg[1] [24]), 
         .Z(key_mem_new_127__N_7264[88])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_51_i89_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_3_lut_4_lut_adj_666 (.A(n33943), .B(n33944), .C(\key_mem_ctrl.num_rounds[2] ), 
         .D(n28850), .Z(clk_c_enable_2413)) /* synthesis lut_function=(A (D)+!A (B (D)+!B !(C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam i1_3_lut_4_lut_adj_666.init = 16'hef00;
    LUT4 mux_51_i80_3_lut_4_lut (.A(n33943), .B(n33944), .C(n33732), .D(\key_reg[1] [15]), 
         .Z(key_mem_new_127__N_7264[79])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_51_i80_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_51_i79_3_lut_4_lut (.A(n33943), .B(n33944), .C(n33733), .D(\key_reg[1] [14]), 
         .Z(key_mem_new_127__N_7264[78])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_51_i79_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_51_i75_3_lut_4_lut (.A(n33943), .B(n33944), .C(n33737), .D(\key_reg[1] [10]), 
         .Z(key_mem_new_127__N_7264[74])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_51_i75_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_51_i67_3_lut_4_lut (.A(n33943), .B(n33944), .C(n33745), .D(\key_reg[1] [2]), 
         .Z(key_mem_new_127__N_7264[66])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_51_i67_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_51_i66_3_lut_4_lut (.A(n33943), .B(n33944), .C(n33746), .D(\key_reg[1] [1]), 
         .Z(key_mem_new_127__N_7264[65])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_51_i66_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25396 (.BLUT(n8_adj_8529), .ALUT(n9_adj_8528), .C0(\muxed_round_nr[1] ), 
          .Z(n30555));
    LUT4 mux_51_i72_3_lut_4_lut (.A(n33943), .B(n33944), .C(n33740), .D(\key_reg[1] [7]), 
         .Z(key_mem_new_127__N_7264[71])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_51_i72_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_51_i83_3_lut_4_lut (.A(n33943), .B(n33944), .C(n33729), .D(\key_reg[1] [18]), 
         .Z(key_mem_new_127__N_7264[82])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_51_i83_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_51_i88_3_lut_4_lut (.A(n33943), .B(n33944), .C(n33724), .D(\key_reg[1] [23]), 
         .Z(key_mem_new_127__N_7264[87])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_51_i88_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_51_i86_3_lut_4_lut (.A(n33943), .B(n33944), .C(n33726), .D(\key_reg[1] [21]), 
         .Z(key_mem_new_127__N_7264[85])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_51_i86_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i35_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [34]), 
         .D(key_mem_new[34]), .Z(key_mem_0__127__N_4960[34])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i35_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_51_i65_3_lut_4_lut (.A(n33943), .B(n33944), .C(n33747), .D(\key_reg[1] [0]), 
         .Z(key_mem_new_127__N_7264[64])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_51_i65_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_51_i68_3_lut_4_lut (.A(n33943), .B(n33944), .C(n33744), .D(\key_reg[1] [3]), 
         .Z(key_mem_new_127__N_7264[67])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_51_i68_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_51_i69_3_lut_4_lut (.A(n33943), .B(n33944), .C(n33743), .D(\key_reg[1] [4]), 
         .Z(key_mem_new_127__N_7264[68])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_51_i69_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_51_i71_3_lut_4_lut (.A(n33943), .B(n33944), .C(n33741), .D(\key_reg[1] [6]), 
         .Z(key_mem_new_127__N_7264[70])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_51_i71_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i10_adj_667 (.BLUT(n2531[3]), .ALUT(n9620), .C0(n29504), .Z(n10_adj_8598));
    LUT4 mux_51_i74_3_lut_4_lut (.A(n33943), .B(n33944), .C(n33738), .D(\key_reg[1] [9]), 
         .Z(key_mem_new_127__N_7264[73])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_51_i74_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_51_i77_3_lut_4_lut (.A(n33943), .B(n33944), .C(n33735), .D(\key_reg[1] [12]), 
         .Z(key_mem_new_127__N_7264[76])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_51_i77_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_51_i127_3_lut_4_lut (.A(n33943), .B(n33944), .C(n33717), 
         .D(\key_reg[0] [30]), .Z(key_mem_new_127__N_7264[126])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_51_i127_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_51_i128_3_lut_4_lut (.A(n33943), .B(n33944), .C(n33716), 
         .D(\key_reg[0] [31]), .Z(key_mem_new_127__N_7264[127])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_51_i128_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_51_i92_3_lut_4_lut (.A(n33943), .B(n33944), .C(n33617), .D(\key_reg[1] [27]), 
         .Z(key_mem_new_127__N_7264[91])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_51_i92_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i1_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [0]), 
         .D(key_mem_new[0]), .Z(key_mem_0__127__N_4960[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i3_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [2]), 
         .D(key_mem_new[2]), .Z(key_mem_0__127__N_4960[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i8_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [7]), 
         .D(key_mem_new[7]), .Z(key_mem_0__127__N_4960[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i7_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [6]), 
         .D(key_mem_new[6]), .Z(key_mem_0__127__N_4960[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i16_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [15]), 
         .D(key_mem_new[15]), .Z(key_mem_0__127__N_4960[15])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i16_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i14_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [13]), 
         .D(key_mem_new[13]), .Z(key_mem_0__127__N_4960[13])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i14_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i20_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [19]), 
         .D(key_mem_new[19]), .Z(key_mem_0__127__N_4960[19])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i20_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i48_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [47]), 
         .D(key_mem_new[47]), .Z(key_mem_0__127__N_4960[47])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i48_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i43_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [42]), 
         .D(key_mem_new[42]), .Z(key_mem_0__127__N_4960[42])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i43_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i53_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [52]), 
         .D(key_mem_new[52]), .Z(key_mem_0__127__N_4960[52])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i53_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25401 (.BLUT(n1_adj_8526), .ALUT(n2_adj_8525), .C0(\muxed_round_nr[1] ), 
          .Z(n30560));
    LUT4 mux_23_i54_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [53]), 
         .D(key_mem_new[53]), .Z(key_mem_0__127__N_4960[53])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i54_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i59_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [58]), 
         .D(key_mem_new[58]), .Z(key_mem_0__127__N_4960[58])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i59_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i64_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [63]), 
         .D(key_mem_new[63]), .Z(key_mem_0__127__N_4960[63])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i64_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i63_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [62]), 
         .D(key_mem_new[62]), .Z(key_mem_0__127__N_4960[62])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i63_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_51_i70_3_lut_4_lut (.A(n33943), .B(n33944), .C(n33742), .D(\key_reg[1] [5]), 
         .Z(key_mem_new_127__N_7264[69])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_51_i70_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_51_i76_3_lut_4_lut (.A(n33943), .B(n33944), .C(n33736), .D(\key_reg[1] [11]), 
         .Z(key_mem_new_127__N_7264[75])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_51_i76_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_51_i78_3_lut_4_lut (.A(n33943), .B(n33944), .C(n33734), .D(\key_reg[1] [13]), 
         .Z(key_mem_new_127__N_7264[77])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_51_i78_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i10_adj_668 (.BLUT(n2531[4]), .ALUT(n9622), .C0(n29504), .Z(n10_adj_8602));
    LUT4 mux_51_i82_3_lut_4_lut (.A(n33943), .B(n33944), .C(n33730), .D(\key_reg[1] [17]), 
         .Z(key_mem_new_127__N_7264[81])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_51_i82_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i13_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [12]), 
         .D(key_mem_new[12]), .Z(key_mem_0__127__N_4960[12])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i13_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25402 (.BLUT(n4_adj_8524), .ALUT(n5_adj_8523), .C0(\muxed_round_nr[1] ), 
          .Z(n30561));
    LUT4 mux_23_i2_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [1]), 
         .D(key_mem_new[1]), .Z(key_mem_0__127__N_4960[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i15_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [14]), 
         .D(key_mem_new[14]), .Z(key_mem_0__127__N_4960[14])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i15_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i17_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [16]), 
         .D(key_mem_new[16]), .Z(key_mem_0__127__N_4960[16])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i17_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i24_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [23]), 
         .D(key_mem_new[23]), .Z(key_mem_0__127__N_4960[23])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i24_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i26_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [25]), 
         .D(key_mem_new[25]), .Z(key_mem_0__127__N_4960[25])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i26_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i25_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [24]), 
         .D(key_mem_new[24]), .Z(key_mem_0__127__N_4960[24])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i25_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i34_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [33]), 
         .D(key_mem_new[33]), .Z(key_mem_0__127__N_4960[33])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i34_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i33_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [32]), 
         .D(key_mem_new[32]), .Z(key_mem_0__127__N_4960[32])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i33_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i40_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [39]), 
         .D(key_mem_new[39]), .Z(key_mem_0__127__N_4960[39])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i40_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_51_i73_3_lut_4_lut (.A(n33943), .B(n33944), .C(n33739), .D(\key_reg[1] [8]), 
         .Z(key_mem_new_127__N_7264[72])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_51_i73_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_51_i87_3_lut_4_lut (.A(n33943), .B(n33944), .C(n33725), .D(\key_reg[1] [22]), 
         .Z(key_mem_new_127__N_7264[86])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_51_i87_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25403 (.BLUT(n8_adj_8522), .ALUT(n9_adj_8521), .C0(\muxed_round_nr[1] ), 
          .Z(n30562));
    LUT4 mux_51_i122_3_lut_4_lut (.A(n33943), .B(n33944), .C(n33722), 
         .D(\key_reg[0] [25]), .Z(key_mem_new_127__N_7264[121])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_51_i122_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i10_adj_669 (.BLUT(n2531[5]), .ALUT(n9624), .C0(n29504), .Z(n10_adj_8607));
    LUT4 mux_23_i5_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [4]), 
         .D(key_mem_new[4]), .Z(key_mem_0__127__N_4960[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i4_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [3]), 
         .D(key_mem_new[3]), .Z(key_mem_0__127__N_4960[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i9_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [8]), 
         .D(key_mem_new[8]), .Z(key_mem_0__127__N_4960[8])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i9_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i6_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [5]), 
         .D(key_mem_new[5]), .Z(key_mem_0__127__N_4960[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i10_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [9]), 
         .D(key_mem_new[9]), .Z(key_mem_0__127__N_4960[9])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i10_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i11_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [10]), 
         .D(key_mem_new[10]), .Z(key_mem_0__127__N_4960[10])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i11_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i18_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [17]), 
         .D(key_mem_new[17]), .Z(key_mem_0__127__N_4960[17])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i18_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i12_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [11]), 
         .D(key_mem_new[11]), .Z(key_mem_0__127__N_4960[11])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i12_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i21_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [20]), 
         .D(key_mem_new[20]), .Z(key_mem_0__127__N_4960[20])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i21_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i19_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [18]), 
         .D(key_mem_new[18]), .Z(key_mem_0__127__N_4960[18])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i19_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i23_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [22]), 
         .D(key_mem_new[22]), .Z(key_mem_0__127__N_4960[22])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i23_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i22_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [21]), 
         .D(key_mem_new[21]), .Z(key_mem_0__127__N_4960[21])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i22_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i27_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [26]), 
         .D(key_mem_new[26]), .Z(key_mem_0__127__N_4960[26])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i27_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i28_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [27]), 
         .D(key_mem_new[27]), .Z(key_mem_0__127__N_4960[27])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i28_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i30_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [29]), 
         .D(key_mem_new[29]), .Z(key_mem_0__127__N_4960[29])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i30_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25408 (.BLUT(n1_adj_8519), .ALUT(n2_adj_8518), .C0(\muxed_round_nr[1] ), 
          .Z(n30567));
    LUT4 mux_23_i29_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [28]), 
         .D(key_mem_new[28]), .Z(key_mem_0__127__N_4960[28])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i29_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i10_adj_670 (.BLUT(n2531[6]), .ALUT(n9626), .C0(n29504), .Z(n10_adj_8608));
    LUT4 mux_23_i32_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [31]), 
         .D(key_mem_new[31]), .Z(key_mem_0__127__N_4960[31])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i32_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i31_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [30]), 
         .D(key_mem_new[30]), .Z(key_mem_0__127__N_4960[30])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i31_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25409 (.BLUT(n4_adj_8517), .ALUT(n5_adj_8516), .C0(\muxed_round_nr[1] ), 
          .Z(n30568));
    LUT4 mux_23_i37_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [36]), 
         .D(key_mem_new[36]), .Z(key_mem_0__127__N_4960[36])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i37_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i36_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [35]), 
         .D(key_mem_new[35]), .Z(key_mem_0__127__N_4960[35])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i36_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i38_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [37]), 
         .D(key_mem_new[37]), .Z(key_mem_0__127__N_4960[37])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i38_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i39_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [38]), 
         .D(key_mem_new[38]), .Z(key_mem_0__127__N_4960[38])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i39_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i42_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [41]), 
         .D(key_mem_new[41]), .Z(key_mem_0__127__N_4960[41])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i42_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i41_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [40]), 
         .D(key_mem_new[40]), .Z(key_mem_0__127__N_4960[40])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i41_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i45_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [44]), 
         .D(key_mem_new[44]), .Z(key_mem_0__127__N_4960[44])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i45_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i44_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [43]), 
         .D(key_mem_new[43]), .Z(key_mem_0__127__N_4960[43])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i44_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i47_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [46]), 
         .D(key_mem_new[46]), .Z(key_mem_0__127__N_4960[46])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i47_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i46_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [45]), 
         .D(key_mem_new[45]), .Z(key_mem_0__127__N_4960[45])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i46_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i10_adj_671 (.BLUT(n2531[7]), .ALUT(n9628), .C0(n29504), .Z(n10_adj_8614));
    LUT4 mux_23_i49_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [48]), 
         .D(key_mem_new[48]), .Z(key_mem_0__127__N_4960[48])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i49_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i50_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [49]), 
         .D(key_mem_new[49]), .Z(key_mem_0__127__N_4960[49])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i50_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i52_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [51]), 
         .D(key_mem_new[51]), .Z(key_mem_0__127__N_4960[51])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i52_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i51_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [50]), 
         .D(key_mem_new[50]), .Z(key_mem_0__127__N_4960[50])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i51_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i56_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [55]), 
         .D(key_mem_new[55]), .Z(key_mem_0__127__N_4960[55])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i56_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i55_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [54]), 
         .D(key_mem_new[54]), .Z(key_mem_0__127__N_4960[54])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i55_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i58_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [57]), 
         .D(key_mem_new[57]), .Z(key_mem_0__127__N_4960[57])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i58_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i57_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [56]), 
         .D(key_mem_new[56]), .Z(key_mem_0__127__N_4960[56])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i57_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i25410 (.BLUT(n8_adj_8515), .ALUT(n9_adj_8514), .C0(\muxed_round_nr[1] ), 
          .Z(n30569));
    LUT4 mux_23_i60_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [59]), 
         .D(key_mem_new[59]), .Z(key_mem_0__127__N_4960[59])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i60_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i61_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [60]), 
         .D(key_mem_new[60]), .Z(key_mem_0__127__N_4960[60])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i61_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i62_3_lut_4_lut (.A(n33943), .B(n33944), .C(\key_mem[0] [61]), 
         .D(key_mem_new[61]), .Z(key_mem_0__127__N_4960[61])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(258[21:39])
    defparam mux_23_i62_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i10_adj_672 (.BLUT(n2531[8]), .ALUT(n9630), .C0(n29504), .Z(n10_adj_8615));
    PFUMX i25415 (.BLUT(n1_adj_8512), .ALUT(n2_adj_8511), .C0(\muxed_round_nr[1] ), 
          .Z(n30574));
    PFUMX i10_adj_673 (.BLUT(n2531[9]), .ALUT(n9632), .C0(n29504), .Z(n10_adj_8617));
    PFUMX i25416 (.BLUT(n4_adj_8510), .ALUT(n5_adj_8509), .C0(\muxed_round_nr[1] ), 
          .Z(n30575));
    LUT4 i14318_2_lut_rep_607 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .Z(n33911)) /* synthesis lut_function=(A (B)) */ ;
    defparam i14318_2_lut_rep_607.init = 16'h8888;
    LUT4 equal_141_i5_2_lut_rep_608 (.A(n35834), .B(round_ctr_reg[1]), .Z(n33912)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam equal_141_i5_2_lut_rep_608.init = 16'hbbbb;
    PFUMX i25417 (.BLUT(n8_adj_8507), .ALUT(n9_adj_8506), .C0(\muxed_round_nr[1] ), 
          .Z(n30576));
    PFUMX i10_adj_674 (.BLUT(n2531[10]), .ALUT(n9634), .C0(n29504), .Z(n10_adj_8620));
    LUT4 mux_85_i88_3_lut_rep_230_4_lut (.A(prev_key0_reg[87]), .B(n4_adj_8421), 
         .C(n33859), .D(\key_reg[5] [23]), .Z(n33534)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam mux_85_i88_3_lut_rep_230_4_lut.init = 16'h6f60;
    LUT4 equal_147_i6_2_lut_rep_612 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .Z(n33916)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam equal_147_i6_2_lut_rep_612.init = 16'hdddd;
    PFUMX i25422 (.BLUT(n1_adj_8504), .ALUT(n2_adj_8503), .C0(\muxed_round_nr[1] ), 
          .Z(n30581));
    PFUMX i10_adj_675 (.BLUT(n2531[11]), .ALUT(n9636), .C0(n29504), .Z(n10_adj_8622));
    PFUMX i25423 (.BLUT(n4_adj_8501), .ALUT(n5_adj_8500), .C0(\muxed_round_nr[1] ), 
          .Z(n30582));
    LUT4 i6_2_lut_3_lut_adj_676 (.A(prev_key1_reg[54]), .B(n33725), .C(keymem_sboxw[22]), 
         .Z(n16677)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;
    defparam i6_2_lut_3_lut_adj_676.init = 16'h9696;
    PFUMX i25424 (.BLUT(n8_adj_8499), .ALUT(n9_adj_8498), .C0(\muxed_round_nr[1] ), 
          .Z(n30583));
    PFUMX i10_adj_677 (.BLUT(n2531[12]), .ALUT(n9638), .C0(n29504), .Z(n10_adj_8625));
    LUT4 i2_2_lut_rep_319 (.A(prev_key0_reg[86]), .B(n4_adj_8417), .Z(n33623)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i2_2_lut_rep_319.init = 16'h6666;
    LUT4 mux_85_i87_3_lut_rep_231_4_lut (.A(prev_key0_reg[86]), .B(n4_adj_8417), 
         .C(n33859), .D(\key_reg[5] [22]), .Z(n33535)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam mux_85_i87_3_lut_rep_231_4_lut.init = 16'h6f60;
    LUT4 i6_2_lut_3_lut_adj_678 (.A(prev_key1_reg[53]), .B(n33726), .C(keymem_sboxw[21]), 
         .Z(n16617)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;
    defparam i6_2_lut_3_lut_adj_678.init = 16'h9696;
    PFUMX i10_adj_679 (.BLUT(n2531[13]), .ALUT(n9640), .C0(n29504), .Z(n10_adj_8627));
    LUT4 i2_2_lut_rep_321 (.A(prev_key0_reg[85]), .B(n4_adj_8410), .Z(n33625)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i2_2_lut_rep_321.init = 16'h6666;
    LUT4 mux_85_i86_3_lut_rep_232_4_lut (.A(prev_key0_reg[85]), .B(n4_adj_8410), 
         .C(n33859), .D(\key_reg[5] [21]), .Z(n33536)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam mux_85_i86_3_lut_rep_232_4_lut.init = 16'h6f60;
    PFUMX i25429 (.BLUT(n1_adj_8496), .ALUT(n2_adj_8495), .C0(\muxed_round_nr[1] ), 
          .Z(n30588));
    PFUMX i25430 (.BLUT(n4_adj_8494), .ALUT(n5_adj_8493), .C0(\muxed_round_nr[1] ), 
          .Z(n30589));
    PFUMX i25431 (.BLUT(n8_adj_8492), .ALUT(n9_adj_8491), .C0(\muxed_round_nr[1] ), 
          .Z(n30590));
    LUT4 i6_2_lut_3_lut_adj_680 (.A(prev_key1_reg[52]), .B(n33727), .C(keymem_sboxw[20]), 
         .Z(n16557)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;
    defparam i6_2_lut_3_lut_adj_680.init = 16'h9696;
    LUT4 i2_2_lut_rep_323 (.A(prev_key0_reg[84]), .B(n4_adj_8403), .Z(n33627)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i2_2_lut_rep_323.init = 16'h6666;
    LUT4 round_3__I_0_Mux_116_i4_3_lut (.A(\key_mem[4] [116]), .B(\key_mem[5] [116]), 
         .C(n33952), .Z(n4_adj_8956)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_116_i4_3_lut.init = 16'hcaca;
    LUT4 mux_85_i85_3_lut_rep_233_4_lut (.A(prev_key0_reg[84]), .B(n4_adj_8403), 
         .C(n33859), .D(\key_reg[5] [20]), .Z(n33537)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam mux_85_i85_3_lut_rep_233_4_lut.init = 16'h6f60;
    PFUMX i25436 (.BLUT(n1_adj_8488), .ALUT(n2_adj_8487), .C0(\muxed_round_nr[1] ), 
          .Z(n30595));
    PFUMX i25437 (.BLUT(n4_adj_8486), .ALUT(n5_adj_8485), .C0(\muxed_round_nr[1] ), 
          .Z(n30596));
    PFUMX i25438 (.BLUT(n8_adj_8484), .ALUT(n9_adj_8483), .C0(\muxed_round_nr[1] ), 
          .Z(n30597));
    LUT4 i6_2_lut_3_lut_adj_681 (.A(prev_key1_reg[51]), .B(n33728), .C(keymem_sboxw[19]), 
         .Z(n16497)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;
    defparam i6_2_lut_3_lut_adj_681.init = 16'h9696;
    LUT4 i15023_2_lut_4_lut (.A(\key_reg[5] [20]), .B(n33627), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[84])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15023_2_lut_4_lut.init = 16'hca00;
    PFUMX i25443 (.BLUT(n1_adj_8481), .ALUT(n2_adj_8480), .C0(\muxed_round_nr[1] ), 
          .Z(n30602));
    PFUMX i25444 (.BLUT(n4_adj_8479), .ALUT(n5_adj_8478), .C0(\muxed_round_nr[1] ), 
          .Z(n30603));
    LUT4 i2_2_lut_rep_325 (.A(prev_key0_reg[83]), .B(n4_adj_8400), .Z(n33629)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i2_2_lut_rep_325.init = 16'h6666;
    LUT4 mux_85_i84_3_lut_rep_234_4_lut (.A(prev_key0_reg[83]), .B(n4_adj_8400), 
         .C(n33859), .D(\key_reg[5] [19]), .Z(n33538)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam mux_85_i84_3_lut_rep_234_4_lut.init = 16'h6f60;
    PFUMX i25445 (.BLUT(n8_adj_8477), .ALUT(n9_adj_8475), .C0(\muxed_round_nr[1] ), 
          .Z(n30604));
    LUT4 i6_2_lut_3_lut_adj_682 (.A(prev_key1_reg[50]), .B(n33729), .C(keymem_sboxw[18]), 
         .Z(n16437)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;
    defparam i6_2_lut_3_lut_adj_682.init = 16'h9696;
    LUT4 i2_2_lut_rep_327 (.A(prev_key0_reg[82]), .B(n4_adj_8395), .Z(n33631)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i2_2_lut_rep_327.init = 16'h6666;
    LUT4 mux_85_i83_3_lut_rep_235_4_lut (.A(prev_key0_reg[82]), .B(n4_adj_8395), 
         .C(n33859), .D(\key_reg[5] [18]), .Z(n33539)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam mux_85_i83_3_lut_rep_235_4_lut.init = 16'h6f60;
    PFUMX i25450 (.BLUT(n1_adj_8470), .ALUT(n2_adj_8469), .C0(\muxed_round_nr[1] ), 
          .Z(n30609));
    PFUMX i25451 (.BLUT(n4_adj_8468), .ALUT(n5_adj_8466), .C0(\muxed_round_nr[1] ), 
          .Z(n30610));
    LUT4 i6_2_lut_3_lut_adj_683 (.A(prev_key1_reg[49]), .B(n33730), .C(keymem_sboxw[17]), 
         .Z(n16377)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;
    defparam i6_2_lut_3_lut_adj_683.init = 16'h9696;
    PFUMX i25452 (.BLUT(n8_adj_8465), .ALUT(n9_adj_8464), .C0(\muxed_round_nr[1] ), 
          .Z(n30611));
    LUT4 i2_2_lut_rep_329 (.A(prev_key0_reg[81]), .B(n4_adj_8390), .Z(n33633)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i2_2_lut_rep_329.init = 16'h6666;
    PFUMX i25457 (.BLUT(n1_adj_8462), .ALUT(n2_adj_8460), .C0(\muxed_round_nr[1] ), 
          .Z(n30616));
    PFUMX i10_adj_684 (.BLUT(n2531[14]), .ALUT(n9642), .C0(n29504), .Z(n10_adj_8633));
    LUT4 equal_140_i6_2_lut_rep_633 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .Z(n33937)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam equal_140_i6_2_lut_rep_633.init = 16'hbbbb;
    PFUMX i10_adj_685 (.BLUT(n2531[15]), .ALUT(n9644), .C0(n29504), .Z(n10_adj_8637));
    LUT4 i14320_2_lut_rep_634 (.A(n35834), .B(round_ctr_reg[1]), .Z(n33938)) /* synthesis lut_function=(A (B)) */ ;
    defparam i14320_2_lut_rep_634.init = 16'h8888;
    PFUMX i25458 (.BLUT(n4_adj_8459), .ALUT(n5_adj_8458), .C0(\muxed_round_nr[1] ), 
          .Z(n30617));
    LUT4 i20116_3_lut_4_lut (.A(round_ctr_reg[0]), .B(round_ctr_reg[1]), 
         .C(round_ctr_reg[2]), .D(round_ctr_reg[3]), .Z(n3[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;
    defparam i20116_3_lut_4_lut.init = 16'h7f80;
    PFUMX i10_adj_686 (.BLUT(n2531[16]), .ALUT(n9646), .C0(n29504), .Z(n10_adj_8639));
    LUT4 i20109_2_lut_3_lut (.A(round_ctr_reg[0]), .B(round_ctr_reg[1]), 
         .C(round_ctr_reg[2]), .Z(n3[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;
    defparam i20109_2_lut_3_lut.init = 16'h7878;
    PFUMX i25459 (.BLUT(n8_adj_8456), .ALUT(n9_adj_8454), .C0(\muxed_round_nr[1] ), 
          .Z(n30618));
    PFUMX i10_adj_687 (.BLUT(n2531[17]), .ALUT(n9648), .C0(n29504), .Z(n10_adj_8640));
    LUT4 mux_85_i82_3_lut_rep_236_4_lut (.A(prev_key0_reg[81]), .B(n4_adj_8390), 
         .C(n33859), .D(\key_reg[5] [17]), .Z(n33540)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam mux_85_i82_3_lut_rep_236_4_lut.init = 16'h6f60;
    LUT4 i6_2_lut_3_lut_adj_688 (.A(prev_key1_reg[48]), .B(n33731), .C(keymem_sboxw[16]), 
         .Z(n16317)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;
    defparam i6_2_lut_3_lut_adj_688.init = 16'h9696;
    LUT4 i2_2_lut_rep_331 (.A(prev_key0_reg[80]), .B(n4_adj_8386), .Z(n33635)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i2_2_lut_rep_331.init = 16'h6666;
    PFUMX i25464 (.BLUT(n1_adj_8452), .ALUT(n2_adj_8450), .C0(\muxed_round_nr[1] ), 
          .Z(n30623));
    LUT4 mux_85_i81_3_lut_rep_237_4_lut (.A(prev_key0_reg[80]), .B(n4_adj_8386), 
         .C(n33859), .D(\key_reg[5] [16]), .Z(n33541)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam mux_85_i81_3_lut_rep_237_4_lut.init = 16'h6f60;
    PFUMX i10_adj_689 (.BLUT(n2531[18]), .ALUT(n9650), .C0(n29504), .Z(n10_adj_8642));
    PFUMX i25465 (.BLUT(n4_adj_8447), .ALUT(n5_adj_8445), .C0(\muxed_round_nr[1] ), 
          .Z(n30624));
    LUT4 equal_147_i5_2_lut_rep_639 (.A(n35834), .B(round_ctr_reg[1]), .Z(n33943)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam equal_147_i5_2_lut_rep_639.init = 16'heeee;
    PFUMX i25605 (.BLUT(n4_adj_8448), .ALUT(n5_adj_8446), .C0(\muxed_round_nr[1] ), 
          .Z(n30764));
    LUT4 i1_2_lut_3_lut_4_lut (.A(n35834), .B(round_ctr_reg[1]), .C(n15483), 
         .D(n33944), .Z(n15484)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_690 (.A(n35834), .B(round_ctr_reg[1]), 
         .C(n15310), .D(n33944), .Z(n15311)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_690.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_691 (.A(n35834), .B(round_ctr_reg[1]), 
         .C(n15423), .D(n33944), .Z(n15424)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_691.init = 16'hf0e0;
    PFUMX i25606 (.BLUT(n8_adj_8443), .ALUT(n9_adj_8442), .C0(\muxed_round_nr[1] ), 
          .Z(n30765));
    LUT4 i1_2_lut_3_lut_4_lut_adj_692 (.A(n35834), .B(round_ctr_reg[1]), 
         .C(n15543), .D(n33944), .Z(n15544)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_692.init = 16'hf0e0;
    LUT4 i6_2_lut_3_lut_adj_693 (.A(prev_key1_reg[47]), .B(n33732), .C(keymem_sboxw[15]), 
         .Z(n16257)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;
    defparam i6_2_lut_3_lut_adj_693.init = 16'h9696;
    LUT4 i1_2_lut_3_lut_4_lut_adj_694 (.A(n35834), .B(round_ctr_reg[1]), 
         .C(n15603), .D(n33944), .Z(n15604)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_694.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_695 (.A(n35834), .B(round_ctr_reg[1]), 
         .C(n15663), .D(n33944), .Z(n15664)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_695.init = 16'hf0e0;
    PFUMX i25466 (.BLUT(n8_adj_8440), .ALUT(n9_adj_8436), .C0(\muxed_round_nr[1] ), 
          .Z(n30625));
    LUT4 i1_2_lut_3_lut_4_lut_adj_696 (.A(n35834), .B(round_ctr_reg[1]), 
         .C(n15723), .D(n33944), .Z(n15724)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_696.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_697 (.A(n35834), .B(round_ctr_reg[1]), 
         .C(n15783), .D(n33944), .Z(n15784)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_697.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_698 (.A(n35834), .B(round_ctr_reg[1]), 
         .C(n15843), .D(n33944), .Z(n15844)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_698.init = 16'hf0e0;
    PFUMX i25611 (.BLUT(n1_adj_8439), .ALUT(n2_adj_8437), .C0(\muxed_round_nr[1] ), 
          .Z(n30770));
    LUT4 i1_2_lut_3_lut_4_lut_adj_699 (.A(n35834), .B(round_ctr_reg[1]), 
         .C(n15903), .D(n33944), .Z(n15904)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_699.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_700 (.A(n35834), .B(round_ctr_reg[1]), 
         .C(n15963), .D(n33944), .Z(n15964)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_700.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_701 (.A(n35834), .B(round_ctr_reg[1]), 
         .C(n16023), .D(n33944), .Z(n16024)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_701.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_702 (.A(n35834), .B(round_ctr_reg[1]), 
         .C(n16083), .D(n33944), .Z(n16084)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_702.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_703 (.A(n35834), .B(round_ctr_reg[1]), 
         .C(n16143), .D(n33944), .Z(n16144)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_703.init = 16'hf0e0;
    PFUMX i25612 (.BLUT(n4_adj_8435), .ALUT(n5_adj_8434), .C0(\muxed_round_nr[1] ), 
          .Z(n30771));
    PFUMX i25613 (.BLUT(n8_adj_8433), .ALUT(n9_adj_8432), .C0(\muxed_round_nr[1] ), 
          .Z(n30772));
    LUT4 i2_2_lut_rep_333 (.A(prev_key0_reg[79]), .B(n4_adj_8381), .Z(n33637)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i2_2_lut_rep_333.init = 16'h6666;
    LUT4 i15022_2_lut_4_lut (.A(\key_reg[5] [19]), .B(n33629), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[83])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15022_2_lut_4_lut.init = 16'hca00;
    PFUMX i25618 (.BLUT(n1_adj_8427), .ALUT(n2_adj_8426), .C0(\muxed_round_nr[1] ), 
          .Z(n30777));
    PFUMX i25471 (.BLUT(n1_adj_8425), .ALUT(n2_adj_8422), .C0(\muxed_round_nr[1] ), 
          .Z(n30630));
    PFUMX i25619 (.BLUT(n4_adj_8424), .ALUT(n5_adj_8423), .C0(\muxed_round_nr[1] ), 
          .Z(n30778));
    PFUMX i25620 (.BLUT(n8_adj_8420), .ALUT(n9_adj_8419), .C0(\muxed_round_nr[1] ), 
          .Z(n30779));
    PFUMX i25472 (.BLUT(n4_adj_8416), .ALUT(n5_adj_8413), .C0(\muxed_round_nr[1] ), 
          .Z(n30631));
    PFUMX i25625 (.BLUT(n1_adj_8415), .ALUT(n2_adj_8414), .C0(\muxed_round_nr[1] ), 
          .Z(n30784));
    PFUMX i25626 (.BLUT(n4_adj_8412), .ALUT(n5_adj_8411), .C0(\muxed_round_nr[1] ), 
          .Z(n30785));
    LUT4 mux_85_i80_3_lut_rep_238_4_lut (.A(prev_key0_reg[79]), .B(n4_adj_8381), 
         .C(n33859), .D(\key_reg[5] [15]), .Z(n33542)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam mux_85_i80_3_lut_rep_238_4_lut.init = 16'h6f60;
    PFUMX i25627 (.BLUT(n8_adj_8408), .ALUT(n9_adj_8407), .C0(\muxed_round_nr[1] ), 
          .Z(n30786));
    PFUMX i25473 (.BLUT(n8_adj_8409), .ALUT(n9_adj_8404), .C0(\muxed_round_nr[1] ), 
          .Z(n30632));
    PFUMX i25632 (.BLUT(n1_adj_8402), .ALUT(n2_adj_8401), .C0(\muxed_round_nr[1] ), 
          .Z(n30791));
    PFUMX i25633 (.BLUT(n4_adj_8399), .ALUT(n5_adj_8398), .C0(\muxed_round_nr[1] ), 
          .Z(n30792));
    PFUMX i25634 (.BLUT(n8_adj_8397), .ALUT(n9_adj_8396), .C0(\muxed_round_nr[1] ), 
          .Z(n30793));
    PFUMX i10_adj_704 (.BLUT(n2531[19]), .ALUT(n9652), .C0(n29504), .Z(n10_adj_8644));
    PFUMX i25639 (.BLUT(n1_adj_8393), .ALUT(n2_adj_8392), .C0(\muxed_round_nr[1] ), 
          .Z(n30798));
    PFUMX i25640 (.BLUT(n4_adj_8389), .ALUT(n5_adj_8388), .C0(\muxed_round_nr[1] ), 
          .Z(n30799));
    LUT4 i6_2_lut_3_lut_adj_705 (.A(prev_key1_reg[46]), .B(n33733), .C(keymem_sboxw[14]), 
         .Z(n16197)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;
    defparam i6_2_lut_3_lut_adj_705.init = 16'h9696;
    PFUMX i25641 (.BLUT(n8_adj_8387), .ALUT(n9_adj_8385), .C0(\muxed_round_nr[1] ), 
          .Z(n30800));
    PFUMX i25646 (.BLUT(n1_adj_8382), .ALUT(n2_adj_8380), .C0(\muxed_round_nr[1] ), 
          .Z(n30805));
    PFUMX i25647 (.BLUT(n4_adj_8379), .ALUT(n5_adj_8378), .C0(\muxed_round_nr[1] ), 
          .Z(n30806));
    PFUMX i25648 (.BLUT(n8_adj_8376), .ALUT(n9_adj_8375), .C0(\muxed_round_nr[1] ), 
          .Z(n30807));
    PFUMX i10_adj_706 (.BLUT(n2531[20]), .ALUT(n9654), .C0(n29504), .Z(n10_adj_8645));
    PFUMX i25478 (.BLUT(n1_adj_8369), .ALUT(n2_adj_8362), .C0(\muxed_round_nr[1] ), 
          .Z(n30637));
    PFUMX i25653 (.BLUT(n1_adj_8372), .ALUT(n2_adj_8371), .C0(\muxed_round_nr[1] ), 
          .Z(n30812));
    PFUMX i25654 (.BLUT(n4_adj_8370), .ALUT(n5_adj_8368), .C0(\muxed_round_nr[1] ), 
          .Z(n30813));
    PFUMX i25655 (.BLUT(n8_adj_8366), .ALUT(n9_adj_8364), .C0(\muxed_round_nr[1] ), 
          .Z(n30814));
    PFUMX i10_adj_707 (.BLUT(n2531[21]), .ALUT(n9656), .C0(n29504), .Z(n10_adj_8648));
    LUT4 i2_2_lut_rep_335 (.A(prev_key0_reg[78]), .B(n4_adj_8377), .Z(n33639)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i2_2_lut_rep_335.init = 16'h6666;
    PFUMX i25660 (.BLUT(n1_adj_8360), .ALUT(n2_adj_8358), .C0(\muxed_round_nr[1] ), 
          .Z(n30819));
    PFUMX i25479 (.BLUT(n4_adj_8354), .ALUT(n5_adj_8351), .C0(\muxed_round_nr[1] ), 
          .Z(n30638));
    PFUMX i25661 (.BLUT(n4_adj_8357), .ALUT(n5_adj_8355), .C0(\muxed_round_nr[1] ), 
          .Z(n30820));
    PFUMX i25662 (.BLUT(n8_adj_8353), .ALUT(n9_adj_8352), .C0(\muxed_round_nr[1] ), 
          .Z(n30821));
    PFUMX i10_adj_708 (.BLUT(n2531[22]), .ALUT(n9658), .C0(n29504), .Z(n10_adj_8650));
    PFUMX i25667 (.BLUT(n1_adj_8345), .ALUT(n2_adj_8344), .C0(\muxed_round_nr[1] ), 
          .Z(n30826));
    PFUMX i25668 (.BLUT(n4_adj_8342), .ALUT(n5_adj_8341), .C0(\muxed_round_nr[1] ), 
          .Z(n30827));
    PFUMX i25480 (.BLUT(n8_adj_8340), .ALUT(n9_adj_8338), .C0(\muxed_round_nr[1] ), 
          .Z(n30639));
    LUT4 i1_2_lut_3_lut_4_lut_adj_709 (.A(n35834), .B(round_ctr_reg[1]), 
         .C(n16203), .D(n33944), .Z(n16204)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_709.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_710 (.A(n35834), .B(round_ctr_reg[1]), 
         .C(n16263), .D(n33944), .Z(n16264)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_710.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_711 (.A(n35834), .B(round_ctr_reg[1]), 
         .C(n16323), .D(n33944), .Z(n16324)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_711.init = 16'hf0e0;
    PFUMX i10_adj_712 (.BLUT(n2531[23]), .ALUT(n9660), .C0(n29504), .Z(n10_adj_8651));
    LUT4 i1_2_lut_3_lut_4_lut_adj_713 (.A(n35834), .B(round_ctr_reg[1]), 
         .C(n16383), .D(n33944), .Z(n16384)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_713.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_714 (.A(n35834), .B(round_ctr_reg[1]), 
         .C(n16443), .D(n33944), .Z(n16444)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_714.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_715 (.A(n35834), .B(round_ctr_reg[1]), 
         .C(n16503), .D(n33944), .Z(n16504)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_715.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_716 (.A(n35834), .B(round_ctr_reg[1]), 
         .C(n16563), .D(n33944), .Z(n16564)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_716.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_717 (.A(n35834), .B(round_ctr_reg[1]), 
         .C(n16623), .D(n33944), .Z(n16624)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_717.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_718 (.A(n35834), .B(round_ctr_reg[1]), 
         .C(n16683), .D(n33944), .Z(n16684)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_718.init = 16'hf0e0;
    PFUMX i25485 (.BLUT(n1_adj_8331), .ALUT(n2_adj_8328), .C0(\muxed_round_nr[1] ), 
          .Z(n30644));
    LUT4 i1_2_lut_3_lut_4_lut_adj_719 (.A(n35834), .B(round_ctr_reg[1]), 
         .C(n16743), .D(n33944), .Z(n16744)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_719.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_720 (.A(n35834), .B(round_ctr_reg[1]), 
         .C(n16803), .D(n33944), .Z(n16804)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_720.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_721 (.A(n35834), .B(round_ctr_reg[1]), 
         .C(n16863), .D(n33944), .Z(n16864)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_721.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_722 (.A(n35834), .B(round_ctr_reg[1]), 
         .C(n16923), .D(n33944), .Z(n16924)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_722.init = 16'hf0e0;
    LUT4 round_3__I_0_Mux_116_i2_3_lut (.A(\key_mem[2] [116]), .B(\key_mem[3] [116]), 
         .C(n33952), .Z(n2_adj_8709)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_116_i2_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_723 (.A(n35834), .B(round_ctr_reg[1]), 
         .C(n16983), .D(n33944), .Z(n16984)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_723.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_724 (.A(n35834), .B(round_ctr_reg[1]), 
         .C(n17043), .D(n33944), .Z(n17044)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_724.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_725 (.A(n35834), .B(round_ctr_reg[1]), 
         .C(n17103), .D(n33944), .Z(n17104)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_725.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_726 (.A(n35834), .B(round_ctr_reg[1]), 
         .C(n17163), .D(n33944), .Z(n17164)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_726.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_727 (.A(n35834), .B(round_ctr_reg[1]), 
         .C(n17223), .D(n33944), .Z(n17224)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_727.init = 16'hf0e0;
    PFUMX i25669 (.BLUT(n8_adj_8330), .ALUT(n9_adj_8329), .C0(\muxed_round_nr[1] ), 
          .Z(n30828));
    PFUMX i10_adj_728 (.BLUT(n2531[24]), .ALUT(n9662), .C0(n29504), .Z(n10_adj_9256));
    LUT4 mux_85_i79_3_lut_rep_239_4_lut (.A(prev_key0_reg[78]), .B(n4_adj_8377), 
         .C(n33859), .D(\key_reg[5] [14]), .Z(n33543)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam mux_85_i79_3_lut_rep_239_4_lut.init = 16'h6f60;
    LUT4 mux_23_i65_4_lut (.A(n35839), .B(\key_mem[0] [64]), .C(n33860), 
         .D(\key_reg[1] [0]), .Z(key_mem_0__127__N_4960[64])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i65_4_lut.init = 16'hcac0;
    PFUMX i25674 (.BLUT(n1_adj_8326), .ALUT(n2_adj_8325), .C0(\muxed_round_nr[1] ), 
          .Z(n30833));
    PFUMX i25486 (.BLUT(n4_adj_8702), .ALUT(n5_adj_8701), .C0(\muxed_round_nr[1] ), 
          .Z(n30645));
    LUT4 mux_23_i66_4_lut (.A(n35839), .B(\key_mem[0] [65]), .C(n33860), 
         .D(\key_reg[1] [1]), .Z(key_mem_0__127__N_4960[65])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i66_4_lut.init = 16'hcac0;
    LUT4 mux_23_i67_4_lut (.A(n35839), .B(\key_mem[0] [66]), .C(n33860), 
         .D(\key_reg[1] [2]), .Z(key_mem_0__127__N_4960[66])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i67_4_lut.init = 16'hcac0;
    LUT4 mux_23_i68_4_lut (.A(n35839), .B(\key_mem[0] [67]), .C(n33860), 
         .D(\key_reg[1] [3]), .Z(key_mem_0__127__N_4960[67])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i68_4_lut.init = 16'hcac0;
    PFUMX i25675 (.BLUT(n4_adj_8324), .ALUT(n5_adj_8323), .C0(\muxed_round_nr[1] ), 
          .Z(n30834));
    LUT4 i1_4_lut_adj_729 (.A(\key_mem_ctrl.num_rounds[2] ), .B(\key_reg[3] [0]), 
         .C(n21_adj_9291), .D(n33860), .Z(prev_key0_new_127__N_4659[0])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(85[17:29])
    defparam i1_4_lut_adj_729.init = 16'ha088;
    LUT4 i6_2_lut_3_lut_adj_730 (.A(prev_key1_reg[45]), .B(n33734), .C(keymem_sboxw[13]), 
         .Z(n16137)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;
    defparam i6_2_lut_3_lut_adj_730.init = 16'h9696;
    LUT4 mux_23_i69_4_lut (.A(n35839), .B(\key_mem[0] [68]), .C(n33860), 
         .D(\key_reg[1] [4]), .Z(key_mem_0__127__N_4960[68])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i69_4_lut.init = 16'hcac0;
    LUT4 mux_23_i70_4_lut (.A(n35839), .B(\key_mem[0] [69]), .C(n33860), 
         .D(\key_reg[1] [5]), .Z(key_mem_0__127__N_4960[69])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i70_4_lut.init = 16'hcac0;
    LUT4 mux_23_i71_4_lut (.A(n35839), .B(\key_mem[0] [70]), .C(n33860), 
         .D(\key_reg[1] [6]), .Z(key_mem_0__127__N_4960[70])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i71_4_lut.init = 16'hcac0;
    PFUMX i25676 (.BLUT(n8_adj_8322), .ALUT(n9_adj_8321), .C0(\muxed_round_nr[1] ), 
          .Z(n30835));
    LUT4 mux_23_i72_4_lut (.A(n35839), .B(\key_mem[0] [71]), .C(n33860), 
         .D(\key_reg[1] [7]), .Z(key_mem_0__127__N_4960[71])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i72_4_lut.init = 16'hcac0;
    LUT4 mux_23_i73_4_lut (.A(n35839), .B(\key_mem[0] [72]), .C(n33860), 
         .D(\key_reg[1] [8]), .Z(key_mem_0__127__N_4960[72])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i73_4_lut.init = 16'hcac0;
    LUT4 mux_23_i74_4_lut (.A(n35839), .B(\key_mem[0] [73]), .C(n33860), 
         .D(\key_reg[1] [9]), .Z(key_mem_0__127__N_4960[73])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i74_4_lut.init = 16'hcac0;
    LUT4 mux_23_i75_4_lut (.A(n35839), .B(\key_mem[0] [74]), .C(n33860), 
         .D(\key_reg[1] [10]), .Z(key_mem_0__127__N_4960[74])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i75_4_lut.init = 16'hcac0;
    LUT4 mux_23_i76_4_lut (.A(n35839), .B(\key_mem[0] [75]), .C(n33860), 
         .D(\key_reg[1] [11]), .Z(key_mem_0__127__N_4960[75])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i76_4_lut.init = 16'hcac0;
    LUT4 i2_2_lut_rep_337 (.A(prev_key0_reg[77]), .B(n4_adj_8373), .Z(n33641)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i2_2_lut_rep_337.init = 16'h6666;
    LUT4 mux_23_i77_4_lut (.A(n35839), .B(\key_mem[0] [76]), .C(n33860), 
         .D(\key_reg[1] [12]), .Z(key_mem_0__127__N_4960[76])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i77_4_lut.init = 16'hcac0;
    LUT4 mux_23_i78_4_lut (.A(n35839), .B(\key_mem[0] [77]), .C(n33860), 
         .D(\key_reg[1] [13]), .Z(key_mem_0__127__N_4960[77])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i78_4_lut.init = 16'hcac0;
    LUT4 mux_23_i79_4_lut (.A(n35839), .B(\key_mem[0] [78]), .C(n33860), 
         .D(\key_reg[1] [14]), .Z(key_mem_0__127__N_4960[78])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i79_4_lut.init = 16'hcac0;
    LUT4 mux_23_i80_4_lut (.A(n35839), .B(\key_mem[0] [79]), .C(n33860), 
         .D(\key_reg[1] [15]), .Z(key_mem_0__127__N_4960[79])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i80_4_lut.init = 16'hcac0;
    LUT4 mux_23_i81_4_lut (.A(n35839), .B(\key_mem[0] [80]), .C(n33860), 
         .D(\key_reg[1] [16]), .Z(key_mem_0__127__N_4960[80])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i81_4_lut.init = 16'hcac0;
    LUT4 mux_23_i82_4_lut (.A(n35839), .B(\key_mem[0] [81]), .C(n33860), 
         .D(\key_reg[1] [17]), .Z(key_mem_0__127__N_4960[81])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i82_4_lut.init = 16'hcac0;
    LUT4 mux_23_i83_4_lut (.A(n35839), .B(\key_mem[0] [82]), .C(n33860), 
         .D(\key_reg[1] [18]), .Z(key_mem_0__127__N_4960[82])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i83_4_lut.init = 16'hcac0;
    LUT4 mux_23_i84_4_lut (.A(n35839), .B(\key_mem[0] [83]), .C(n33860), 
         .D(\key_reg[1] [19]), .Z(key_mem_0__127__N_4960[83])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i84_4_lut.init = 16'hcac0;
    LUT4 mux_23_i85_4_lut (.A(n35839), .B(\key_mem[0] [84]), .C(n33860), 
         .D(\key_reg[1] [20]), .Z(key_mem_0__127__N_4960[84])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i85_4_lut.init = 16'hcac0;
    LUT4 mux_23_i86_4_lut (.A(n35839), .B(\key_mem[0] [85]), .C(n33860), 
         .D(\key_reg[1] [21]), .Z(key_mem_0__127__N_4960[85])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i86_4_lut.init = 16'hcac0;
    LUT4 mux_23_i87_4_lut (.A(n35839), .B(\key_mem[0] [86]), .C(n33860), 
         .D(\key_reg[1] [22]), .Z(key_mem_0__127__N_4960[86])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i87_4_lut.init = 16'hcac0;
    LUT4 mux_23_i88_4_lut (.A(n35839), .B(\key_mem[0] [87]), .C(n33860), 
         .D(\key_reg[1] [23]), .Z(key_mem_0__127__N_4960[87])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i88_4_lut.init = 16'hcac0;
    LUT4 mux_85_i78_3_lut_rep_240_4_lut (.A(prev_key0_reg[77]), .B(n4_adj_8373), 
         .C(n33859), .D(\key_reg[5] [13]), .Z(n33544)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam mux_85_i78_3_lut_rep_240_4_lut.init = 16'h6f60;
    LUT4 i6_2_lut_3_lut_adj_731 (.A(prev_key1_reg[44]), .B(n33735), .C(keymem_sboxw[12]), 
         .Z(n16077)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;
    defparam i6_2_lut_3_lut_adj_731.init = 16'h9696;
    LUT4 equal_148_i6_2_lut_rep_640 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .Z(n33944)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam equal_148_i6_2_lut_rep_640.init = 16'heeee;
    LUT4 i2_2_lut_rep_339 (.A(prev_key0_reg[76]), .B(n4_adj_8367), .Z(n33643)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i2_2_lut_rep_339.init = 16'h6666;
    LUT4 mux_23_i89_4_lut (.A(n35839), .B(\key_mem[0] [88]), .C(n33860), 
         .D(\key_reg[1] [24]), .Z(key_mem_0__127__N_4960[88])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i89_4_lut.init = 16'hcac0;
    LUT4 mux_23_i90_4_lut (.A(n35839), .B(\key_mem[0] [89]), .C(n33860), 
         .D(\key_reg[1] [25]), .Z(key_mem_0__127__N_4960[89])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i90_4_lut.init = 16'hcac0;
    LUT4 mux_23_i91_4_lut (.A(n35839), .B(\key_mem[0] [90]), .C(n33860), 
         .D(\key_reg[1] [26]), .Z(key_mem_0__127__N_4960[90])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i91_4_lut.init = 16'hcac0;
    LUT4 equal_120_i7_2_lut_rep_556_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(round_ctr_reg[1]), .D(n35834), .Z(n33860)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam equal_120_i7_2_lut_rep_556_3_lut_4_lut.init = 16'hfffe;
    LUT4 mux_23_i92_4_lut (.A(n35839), .B(\key_mem[0] [91]), .C(n33860), 
         .D(\key_reg[1] [27]), .Z(key_mem_0__127__N_4960[91])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i92_4_lut.init = 16'hcac0;
    LUT4 mux_23_i93_4_lut (.A(n35839), .B(\key_mem[0] [92]), .C(n33860), 
         .D(\key_reg[1] [28]), .Z(key_mem_0__127__N_4960[92])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i93_4_lut.init = 16'hcac0;
    LUT4 mux_23_i94_4_lut (.A(n35839), .B(\key_mem[0] [93]), .C(n33860), 
         .D(\key_reg[1] [29]), .Z(key_mem_0__127__N_4960[93])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i94_4_lut.init = 16'hcac0;
    LUT4 mux_23_i95_4_lut (.A(n35839), .B(\key_mem[0] [94]), .C(n33860), 
         .D(\key_reg[1] [30]), .Z(key_mem_0__127__N_4960[94])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i95_4_lut.init = 16'hcac0;
    LUT4 mux_23_i96_4_lut (.A(n35839), .B(\key_mem[0] [95]), .C(n33860), 
         .D(\key_reg[1] [31]), .Z(key_mem_0__127__N_4960[95])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i96_4_lut.init = 16'hcac0;
    LUT4 mux_23_i97_4_lut (.A(n35839), .B(\key_mem[0] [96]), .C(n33860), 
         .D(\key_reg[0] [0]), .Z(key_mem_0__127__N_4960[96])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i97_4_lut.init = 16'hcac0;
    LUT4 mux_23_i98_4_lut (.A(n35839), .B(\key_mem[0] [97]), .C(n33860), 
         .D(\key_reg[0] [1]), .Z(key_mem_0__127__N_4960[97])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i98_4_lut.init = 16'hcac0;
    LUT4 mux_23_i99_4_lut (.A(n35839), .B(\key_mem[0] [98]), .C(n33860), 
         .D(\key_reg[0] [2]), .Z(key_mem_0__127__N_4960[98])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i99_4_lut.init = 16'hcac0;
    LUT4 mux_23_i100_4_lut (.A(n35839), .B(\key_mem[0] [99]), .C(n33860), 
         .D(\key_reg[0] [3]), .Z(key_mem_0__127__N_4960[99])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i100_4_lut.init = 16'hcac0;
    LUT4 mux_23_i101_4_lut (.A(n35839), .B(\key_mem[0] [100]), .C(n33860), 
         .D(\key_reg[0] [4]), .Z(key_mem_0__127__N_4960[100])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i101_4_lut.init = 16'hcac0;
    LUT4 mux_23_i102_4_lut (.A(n35839), .B(\key_mem[0] [101]), .C(n33860), 
         .D(\key_reg[0] [5]), .Z(key_mem_0__127__N_4960[101])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i102_4_lut.init = 16'hcac0;
    LUT4 round_3__I_0_Mux_105_i1_3_lut (.A(\key_mem[0] [105]), .B(\key_mem[1] [105]), 
         .C(n33952), .Z(n1)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_105_i1_3_lut.init = 16'hcaca;
    LUT4 mux_23_i103_4_lut (.A(n35839), .B(\key_mem[0] [102]), .C(n33860), 
         .D(\key_reg[0] [6]), .Z(key_mem_0__127__N_4960[102])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i103_4_lut.init = 16'hcac0;
    LUT4 mux_23_i104_4_lut (.A(n35839), .B(\key_mem[0] [103]), .C(n33860), 
         .D(\key_reg[0] [7]), .Z(key_mem_0__127__N_4960[103])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i104_4_lut.init = 16'hcac0;
    LUT4 mux_23_i105_4_lut (.A(n35839), .B(\key_mem[0] [104]), .C(n33860), 
         .D(\key_reg[0] [8]), .Z(key_mem_0__127__N_4960[104])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i105_4_lut.init = 16'hcac0;
    LUT4 mux_23_i106_4_lut (.A(n35839), .B(\key_mem[0] [105]), .C(n33860), 
         .D(\key_reg[0] [9]), .Z(key_mem_0__127__N_4960[105])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i106_4_lut.init = 16'hcac0;
    LUT4 mux_23_i107_4_lut (.A(n35839), .B(\key_mem[0] [106]), .C(n33860), 
         .D(\key_reg[0] [10]), .Z(key_mem_0__127__N_4960[106])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i107_4_lut.init = 16'hcac0;
    LUT4 mux_23_i108_4_lut (.A(n35839), .B(\key_mem[0] [107]), .C(n33860), 
         .D(\key_reg[0] [11]), .Z(key_mem_0__127__N_4960[107])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i108_4_lut.init = 16'hcac0;
    LUT4 mux_23_i109_4_lut (.A(n35839), .B(\key_mem[0] [108]), .C(n33860), 
         .D(\key_reg[0] [12]), .Z(key_mem_0__127__N_4960[108])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i109_4_lut.init = 16'hcac0;
    LUT4 mux_23_i110_4_lut (.A(n35839), .B(\key_mem[0] [109]), .C(n33860), 
         .D(\key_reg[0] [13]), .Z(key_mem_0__127__N_4960[109])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i110_4_lut.init = 16'hcac0;
    LUT4 mux_23_i111_4_lut (.A(n35839), .B(\key_mem[0] [110]), .C(n33860), 
         .D(\key_reg[0] [14]), .Z(key_mem_0__127__N_4960[110])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i111_4_lut.init = 16'hcac0;
    LUT4 mux_23_i112_4_lut (.A(n35839), .B(\key_mem[0] [111]), .C(n33860), 
         .D(\key_reg[0] [15]), .Z(key_mem_0__127__N_4960[111])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i112_4_lut.init = 16'hcac0;
    LUT4 mux_23_i113_4_lut (.A(n35839), .B(\key_mem[0] [112]), .C(n33860), 
         .D(\key_reg[0] [16]), .Z(key_mem_0__127__N_4960[112])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i113_4_lut.init = 16'hcac0;
    LUT4 mux_23_i114_4_lut (.A(n35839), .B(\key_mem[0] [113]), .C(n33860), 
         .D(\key_reg[0] [17]), .Z(key_mem_0__127__N_4960[113])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i114_4_lut.init = 16'hcac0;
    LUT4 mux_23_i115_4_lut (.A(n35839), .B(\key_mem[0] [114]), .C(n33860), 
         .D(\key_reg[0] [18]), .Z(key_mem_0__127__N_4960[114])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i115_4_lut.init = 16'hcac0;
    LUT4 mux_23_i116_4_lut (.A(n35839), .B(\key_mem[0] [115]), .C(n33860), 
         .D(\key_reg[0] [19]), .Z(key_mem_0__127__N_4960[115])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i116_4_lut.init = 16'hcac0;
    LUT4 mux_23_i117_4_lut (.A(n35839), .B(\key_mem[0] [116]), .C(n33860), 
         .D(\key_reg[0] [20]), .Z(key_mem_0__127__N_4960[116])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i117_4_lut.init = 16'hcac0;
    LUT4 mux_23_i118_4_lut (.A(n35839), .B(\key_mem[0] [117]), .C(n33860), 
         .D(\key_reg[0] [21]), .Z(key_mem_0__127__N_4960[117])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i118_4_lut.init = 16'hcac0;
    LUT4 mux_23_i119_4_lut (.A(n35839), .B(\key_mem[0] [118]), .C(n33860), 
         .D(\key_reg[0] [22]), .Z(key_mem_0__127__N_4960[118])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i119_4_lut.init = 16'hcac0;
    LUT4 mux_23_i120_4_lut (.A(n35839), .B(\key_mem[0] [119]), .C(n33860), 
         .D(\key_reg[0] [23]), .Z(key_mem_0__127__N_4960[119])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i120_4_lut.init = 16'hcac0;
    LUT4 mux_23_i121_4_lut (.A(n35839), .B(\key_mem[0] [120]), .C(n33860), 
         .D(\key_reg[0] [24]), .Z(key_mem_0__127__N_4960[120])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i121_4_lut.init = 16'hcac0;
    LUT4 mux_23_i122_4_lut (.A(n35839), .B(\key_mem[0] [121]), .C(n33860), 
         .D(\key_reg[0] [25]), .Z(key_mem_0__127__N_4960[121])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i122_4_lut.init = 16'hcac0;
    LUT4 mux_23_i123_4_lut (.A(n35839), .B(\key_mem[0] [122]), .C(n33860), 
         .D(\key_reg[0] [26]), .Z(key_mem_0__127__N_4960[122])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i123_4_lut.init = 16'hcac0;
    LUT4 mux_23_i124_4_lut (.A(n35839), .B(\key_mem[0] [123]), .C(n33860), 
         .D(\key_reg[0] [27]), .Z(key_mem_0__127__N_4960[123])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i124_4_lut.init = 16'hcac0;
    LUT4 mux_23_i125_4_lut (.A(n35839), .B(\key_mem[0] [124]), .C(n33860), 
         .D(\key_reg[0] [28]), .Z(key_mem_0__127__N_4960[124])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i125_4_lut.init = 16'hcac0;
    LUT4 mux_23_i126_4_lut (.A(n35839), .B(\key_mem[0] [125]), .C(n33860), 
         .D(\key_reg[0] [29]), .Z(key_mem_0__127__N_4960[125])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i126_4_lut.init = 16'hcac0;
    LUT4 mux_23_i127_4_lut (.A(n35839), .B(\key_mem[0] [126]), .C(n33860), 
         .D(\key_reg[0] [30]), .Z(key_mem_0__127__N_4960[126])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i127_4_lut.init = 16'hcac0;
    LUT4 mux_23_i128_4_lut (.A(n35839), .B(\key_mem[0] [127]), .C(n33860), 
         .D(\key_reg[0] [31]), .Z(key_mem_0__127__N_4960[127])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:20])
    defparam mux_23_i128_4_lut.init = 16'hcac0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_732 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[38]), .D(n33945), .Z(n22_adj_8270)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_732.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_733 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[37]), .D(n33945), .Z(n22_adj_8269)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_733.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_734 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[36]), .D(n33945), .Z(n22_adj_8268)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_734.init = 16'hf0e0;
    LUT4 i14997_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[119]), .D(n33945), .Z(n8680[119])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14997_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i14992_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[114]), .D(n33945), .Z(n8680[114])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14992_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i14988_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[110]), .D(n33945), .Z(n8680[110])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14988_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i14324_2_lut (.A(n35839), .B(n6361[2]), .Z(round_ctr_we)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(350[12] 354[12])
    defparam i14324_2_lut.init = 16'heeee;
    LUT4 i20102_2_lut (.A(round_ctr_reg[1]), .B(round_ctr_reg[0]), .Z(n3[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(352[27:47])
    defparam i20102_2_lut.init = 16'h6666;
    LUT4 round_3__I_0_Mux_104_i11_3_lut (.A(\key_mem[12] [104]), .B(\key_mem[13] [104]), 
         .C(n33952), .Z(n11_adj_127)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_104_i11_3_lut.init = 16'hcaca;
    LUT4 round_3__I_0_Mux_104_i9_3_lut (.A(\key_mem[10] [104]), .B(\key_mem[11] [104]), 
         .C(n33952), .Z(n9)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_104_i9_3_lut.init = 16'hcaca;
    LUT4 i14983_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[105]), .D(n33945), .Z(n8680[105])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14983_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i9476_1_lut (.A(n35839), .Z(n15086)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam i9476_1_lut.init = 16'h5555;
    LUT4 rcon_reg_6__I_0_i5_2_lut (.A(rcon_reg[3]), .B(\rcon_logic.tmp_rcon [0]), 
         .Z(\rcon_logic.tmp_rcon [4])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(318[18:70])
    defparam rcon_reg_6__I_0_i5_2_lut.init = 16'h6666;
    LUT4 rcon_reg_6__I_0_i2_2_lut (.A(rcon_reg[0]), .B(\rcon_logic.tmp_rcon [0]), 
         .Z(\rcon_logic.tmp_rcon [1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(318[18:70])
    defparam rcon_reg_6__I_0_i2_2_lut.init = 16'h6666;
    LUT4 i1074_1_lut (.A(round_ctr_reg[0]), .Z(n1_adj_9290)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1074_1_lut.init = 16'h5555;
    LUT4 i1_2_lut_adj_735 (.A(prev_key0_reg[24]), .B(prev_key0_reg[56]), 
         .Z(n4_adj_9084)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_adj_735.init = 16'h6666;
    LUT4 i1_2_lut_adj_736 (.A(prev_key0_reg[25]), .B(prev_key0_reg[57]), 
         .Z(n4_adj_9067)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_adj_736.init = 16'h6666;
    LUT4 i1_2_lut_adj_737 (.A(prev_key0_reg[26]), .B(prev_key0_reg[58]), 
         .Z(n4_adj_9064)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_adj_737.init = 16'h6666;
    LUT4 i1_2_lut_adj_738 (.A(prev_key0_reg[27]), .B(prev_key0_reg[59]), 
         .Z(n4_adj_9061)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_adj_738.init = 16'h6666;
    LUT4 i14974_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[96]), .D(n33945), .Z(n8680[96])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14974_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i14968_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[90]), .D(n33945), .Z(n8680[90])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14968_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i14964_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[86]), .D(n33945), .Z(n8680[86])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14964_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i1_2_lut_adj_739 (.A(prev_key0_reg[28]), .B(prev_key0_reg[60]), 
         .Z(n4_adj_9059)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_adj_739.init = 16'h6666;
    LUT4 i14960_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[82]), .D(n33945), .Z(n8680[82])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14960_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 round_3__I_0_Mux_104_i8_3_lut (.A(\key_mem[8] [104]), .B(\key_mem[9] [104]), 
         .C(n33952), .Z(n8)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_104_i8_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_740 (.A(prev_key0_reg[29]), .B(prev_key0_reg[61]), 
         .Z(n4_adj_9055)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_adj_740.init = 16'h6666;
    LUT4 i1_2_lut_3_lut_4_lut_adj_741 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(keymem_sboxw[31]), .D(n33945), .Z(n21_adj_8264)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_741.init = 16'hf0e0;
    LUT4 i1_2_lut_adj_742 (.A(prev_key0_reg[30]), .B(prev_key0_reg[62]), 
         .Z(n4_adj_9054)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_adj_742.init = 16'h6666;
    LUT4 i15001_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[124]), .D(n33945), .Z(n8680[124])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i15001_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i14995_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[117]), .D(n33945), .Z(n8680[117])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14995_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i14986_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[108]), .D(n33945), .Z(n8680[108])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14986_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i14981_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[103]), .D(n33945), .Z(n8680[103])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14981_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i1_2_lut_adj_743 (.A(prev_key0_reg[31]), .B(prev_key0_reg[63]), 
         .Z(n4_adj_9051)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_adj_743.init = 16'h6666;
    LUT4 i14979_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[101]), .D(n33945), .Z(n8680[101])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14979_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i14976_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[98]), .D(n33945), .Z(n8680[98])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14976_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i14972_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[94]), .D(n33945), .Z(n8680[94])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14972_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i14969_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[91]), .D(n33945), .Z(n8680[91])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14969_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i14967_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[89]), .D(n33945), .Z(n8680[89])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14967_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i14963_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[85]), .D(n33945), .Z(n8680[85])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14963_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i14959_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[81]), .D(n33945), .Z(n8680[81])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14959_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i1_2_lut_adj_744 (.A(prev_key0_reg[0]), .B(prev_key0_reg[32]), 
         .Z(n4_adj_9048)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_adj_744.init = 16'h6666;
    LUT4 i1_2_lut_3_lut_4_lut_adj_745 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[40]), .D(n33945), .Z(n22_adj_8272)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_745.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_746 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[32]), .D(n33945), .Z(n22)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_746.init = 16'hf0e0;
    LUT4 i14998_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[120]), .D(n33945), .Z(n8680[120])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14998_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i1_2_lut_adj_747 (.A(prev_key0_reg[1]), .B(prev_key0_reg[33]), 
         .Z(n4_adj_9046)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_adj_747.init = 16'h6666;
    LUT4 i14990_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[112]), .D(n33945), .Z(n8680[112])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14990_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i14984_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[106]), .D(n33945), .Z(n8680[106])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14984_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i1_2_lut_adj_748 (.A(prev_key0_reg[2]), .B(prev_key0_reg[34]), 
         .Z(n4_adj_9042)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_adj_748.init = 16'h6666;
    LUT4 i14996_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[118]), .D(n33945), .Z(n8680[118])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14996_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i1_2_lut_adj_749 (.A(prev_key0_reg[3]), .B(prev_key0_reg[35]), 
         .Z(n4_adj_9040)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_adj_749.init = 16'h6666;
    LUT4 i1_2_lut_adj_750 (.A(prev_key0_reg[4]), .B(prev_key0_reg[36]), 
         .Z(n4_adj_9034)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_adj_750.init = 16'h6666;
    LUT4 i1_2_lut_3_lut_4_lut_adj_751 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[54]), .D(n33945), .Z(n22_adj_8286)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_751.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_752 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[53]), .D(n33945), .Z(n22_adj_8285)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_752.init = 16'hf0e0;
    LUT4 i1_2_lut_adj_753 (.A(prev_key0_reg[5]), .B(prev_key0_reg[37]), 
         .Z(n4_adj_9032)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_adj_753.init = 16'h6666;
    LUT4 i1_2_lut_3_lut_4_lut_adj_754 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[52]), .D(n33945), .Z(n22_adj_8284)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_754.init = 16'hf0e0;
    LUT4 i1_2_lut_adj_755 (.A(prev_key0_reg[6]), .B(prev_key0_reg[38]), 
         .Z(n4_adj_9029)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_adj_755.init = 16'h6666;
    LUT4 i1_2_lut_adj_756 (.A(prev_key0_reg[7]), .B(prev_key0_reg[39]), 
         .Z(n4_adj_9027)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_adj_756.init = 16'h6666;
    LUT4 i1_2_lut_3_lut_4_lut_adj_757 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[51]), .D(n33945), .Z(n22_adj_8283)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_757.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_758 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[50]), .D(n33945), .Z(n22_adj_8282)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_758.init = 16'hf0e0;
    LUT4 i1_2_lut_adj_759 (.A(prev_key0_reg[8]), .B(prev_key0_reg[40]), 
         .Z(n4_adj_9024)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_adj_759.init = 16'h6666;
    LUT4 i1_2_lut_3_lut_4_lut_adj_760 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[49]), .D(n33945), .Z(n22_adj_8281)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_760.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_761 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[48]), .D(n33945), .Z(n22_adj_8280)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_761.init = 16'hf0e0;
    LUT4 i1_2_lut_adj_762 (.A(prev_key0_reg[9]), .B(prev_key0_reg[41]), 
         .Z(n4_adj_9021)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_adj_762.init = 16'h6666;
    LUT4 i1_2_lut_3_lut_4_lut_adj_763 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[47]), .D(n33945), .Z(n22_adj_8279)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_763.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_764 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[46]), .D(n33945), .Z(n22_adj_8278)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_764.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_765 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[45]), .D(n33945), .Z(n22_adj_8277)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_765.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_766 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[44]), .D(n33945), .Z(n22_adj_8276)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_766.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_767 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[43]), .D(n33945), .Z(n22_adj_8275)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_767.init = 16'hf0e0;
    LUT4 i1_2_lut_adj_768 (.A(prev_key0_reg[10]), .B(prev_key0_reg[42]), 
         .Z(n4_adj_9019)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_adj_768.init = 16'h6666;
    LUT4 i1_2_lut_adj_769 (.A(prev_key0_reg[11]), .B(prev_key0_reg[43]), 
         .Z(n4_adj_9015)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_adj_769.init = 16'h6666;
    LUT4 i1_2_lut_adj_770 (.A(prev_key0_reg[12]), .B(prev_key0_reg[44]), 
         .Z(n4_adj_9013)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_adj_770.init = 16'h6666;
    LUT4 i1_2_lut_adj_771 (.A(prev_key0_reg[13]), .B(prev_key0_reg[45]), 
         .Z(n4_adj_9011)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_adj_771.init = 16'h6666;
    LUT4 i1_2_lut_adj_772 (.A(prev_key0_reg[14]), .B(prev_key0_reg[46]), 
         .Z(n4_adj_9007)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_adj_772.init = 16'h6666;
    LUT4 i1_2_lut_adj_773 (.A(prev_key0_reg[15]), .B(prev_key0_reg[47]), 
         .Z(n4_adj_9003)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_adj_773.init = 16'h6666;
    LUT4 i1_2_lut_adj_774 (.A(prev_key0_reg[16]), .B(prev_key0_reg[48]), 
         .Z(n4_adj_9001)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_adj_774.init = 16'h6666;
    LUT4 i1_2_lut_adj_775 (.A(prev_key0_reg[17]), .B(prev_key0_reg[49]), 
         .Z(n4_adj_9000)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_adj_775.init = 16'h6666;
    LUT4 i1_2_lut_adj_776 (.A(prev_key0_reg[18]), .B(prev_key0_reg[50]), 
         .Z(n4_adj_8995)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_adj_776.init = 16'h6666;
    LUT4 i1_2_lut_3_lut_4_lut_adj_777 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[42]), .D(n33945), .Z(n22_adj_8274)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_777.init = 16'hf0e0;
    LUT4 i1_2_lut_adj_778 (.A(prev_key0_reg[19]), .B(prev_key0_reg[51]), 
         .Z(n4_adj_8993)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_adj_778.init = 16'h6666;
    LUT4 i1_2_lut_adj_779 (.A(prev_key0_reg[20]), .B(prev_key0_reg[52]), 
         .Z(n4_adj_8990)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_adj_779.init = 16'h6666;
    LUT4 i1_2_lut_3_lut_4_lut_adj_780 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[41]), .D(n33945), .Z(n22_adj_8273)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_780.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_781 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[39]), .D(n33945), .Z(n22_adj_8271)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_781.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_782 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[35]), .D(n33945), .Z(n22_adj_8267)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_782.init = 16'hf0e0;
    LUT4 i1_2_lut_adj_783 (.A(prev_key0_reg[21]), .B(prev_key0_reg[53]), 
         .Z(n4_adj_8988)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_adj_783.init = 16'h6666;
    LUT4 i1_2_lut_adj_784 (.A(prev_key0_reg[22]), .B(prev_key0_reg[54]), 
         .Z(n4_adj_8984)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_adj_784.init = 16'h6666;
    LUT4 i1_2_lut_adj_785 (.A(prev_key0_reg[23]), .B(prev_key0_reg[55]), 
         .Z(n4_adj_8980)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_adj_785.init = 16'h6666;
    LUT4 i1_2_lut_3_lut_4_lut_adj_786 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[34]), .D(n33945), .Z(n22_adj_8266)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_786.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_787 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[33]), .D(n33945), .Z(n22_adj_8265)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_787.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_788 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(keymem_sboxw[30]), .D(n33945), .Z(n21_adj_8263)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_788.init = 16'hf0e0;
    FD1P3AX key_mem_ctrl_reg_FSM_i0_i1_rep_692 (.D(n6361[2]), .SP(key_mem_ctrl_we), 
            .CK(clk_c), .Q(clk_c_enable_2286));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam key_mem_ctrl_reg_FSM_i0_i1_rep_692.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_4_lut_adj_789 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[57]), .D(n33945), .Z(n22_adj_8289)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_789.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_790 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[56]), .D(n33945), .Z(n22_adj_8288)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_790.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_791 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[55]), .D(n33945), .Z(n22_adj_8287)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_791.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_792 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(keymem_sboxw[0]), .D(n33945), .Z(n21_adj_9291)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_792.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_793 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(keymem_sboxw[1]), .D(n33945), .Z(n21)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_793.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_794 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(keymem_sboxw[2]), .D(n33945), .Z(n21_adj_8235)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_794.init = 16'hf0e0;
    FD1P3AX key_mem_ctrl_reg_FSM_i0_i1_rep_691 (.D(n6361[2]), .SP(key_mem_ctrl_we), 
            .CK(clk_c), .Q(clk_c_enable_2236));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam key_mem_ctrl_reg_FSM_i0_i1_rep_691.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_4_lut_adj_795 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(keymem_sboxw[3]), .D(n33945), .Z(n21_adj_8236)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_795.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_796 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(keymem_sboxw[4]), .D(n33945), .Z(n21_adj_8237)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_796.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_797 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(keymem_sboxw[5]), .D(n33945), .Z(n21_adj_8238)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_797.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_798 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(keymem_sboxw[6]), .D(n33945), .Z(n21_adj_8239)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_798.init = 16'hf0e0;
    FD1P3AX key_mem_ctrl_reg_FSM_i0_i1_rep_690 (.D(n6361[2]), .SP(key_mem_ctrl_we), 
            .CK(clk_c), .Q(clk_c_enable_2186));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam key_mem_ctrl_reg_FSM_i0_i1_rep_690.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_4_lut_adj_799 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(keymem_sboxw[7]), .D(n33945), .Z(n21_adj_8240)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_799.init = 16'hf0e0;
    FD1P3AX key_mem_ctrl_reg_FSM_i0_i1_rep_689 (.D(n6361[2]), .SP(key_mem_ctrl_we), 
            .CK(clk_c), .Q(clk_c_enable_2136));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam key_mem_ctrl_reg_FSM_i0_i1_rep_689.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_4_lut_adj_800 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(keymem_sboxw[8]), .D(n33945), .Z(n21_adj_8241)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_800.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_801 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(keymem_sboxw[9]), .D(n33945), .Z(n21_adj_8242)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_801.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_802 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(keymem_sboxw[10]), .D(n33945), .Z(n21_adj_8243)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_802.init = 16'hf0e0;
    FD1P3AX key_mem_ctrl_reg_FSM_i0_i1_rep_688 (.D(n6361[2]), .SP(key_mem_ctrl_we), 
            .CK(clk_c), .Q(clk_c_enable_2086));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam key_mem_ctrl_reg_FSM_i0_i1_rep_688.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_4_lut_adj_803 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(keymem_sboxw[11]), .D(n33945), .Z(n21_adj_8244)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_803.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_804 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(keymem_sboxw[12]), .D(n33945), .Z(n21_adj_8245)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_804.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_805 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(keymem_sboxw[13]), .D(n33945), .Z(n21_adj_8246)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_805.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_806 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(keymem_sboxw[14]), .D(n33945), .Z(n21_adj_8247)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_806.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_807 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(keymem_sboxw[15]), .D(n33945), .Z(n21_adj_8248)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_807.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_808 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(keymem_sboxw[16]), .D(n33945), .Z(n21_adj_8249)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_808.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_809 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(keymem_sboxw[17]), .D(n33945), .Z(n21_adj_8250)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_809.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_810 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(keymem_sboxw[18]), .D(n33945), .Z(n21_adj_8251)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_810.init = 16'hf0e0;
    FD1P3AX key_mem_ctrl_reg_FSM_i0_i1_rep_687 (.D(n6361[2]), .SP(key_mem_ctrl_we), 
            .CK(clk_c), .Q(clk_c_enable_2036));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam key_mem_ctrl_reg_FSM_i0_i1_rep_687.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_4_lut_adj_811 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(keymem_sboxw[19]), .D(n33945), .Z(n21_adj_8252)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_811.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_812 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(keymem_sboxw[20]), .D(n33945), .Z(n21_adj_8253)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_812.init = 16'hf0e0;
    PFUMX i10_adj_813 (.BLUT(n2531[25]), .ALUT(n9664), .C0(n29504), .Z(n10_adj_9258));
    LUT4 i1_2_lut_3_lut_4_lut_adj_814 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(keymem_sboxw[21]), .D(n33945), .Z(n21_adj_8254)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_814.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_815 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(keymem_sboxw[22]), .D(n33945), .Z(n21_adj_8255)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_815.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_816 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(keymem_sboxw[23]), .D(n33945), .Z(n21_adj_8256)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_816.init = 16'hf0e0;
    FD1P3AX key_mem_ctrl_reg_FSM_i0_i1_rep_686 (.D(n6361[2]), .SP(key_mem_ctrl_we), 
            .CK(clk_c), .Q(clk_c_enable_1986));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam key_mem_ctrl_reg_FSM_i0_i1_rep_686.GSR = "ENABLED";
    PFUMX i25487 (.BLUT(n8_adj_8700), .ALUT(n9_adj_8699), .C0(\muxed_round_nr[1] ), 
          .Z(n30646));
    PFUMX i10_adj_817 (.BLUT(n2531[26]), .ALUT(n9666), .C0(n29504), .Z(n10_adj_9260));
    PFUMX i10_adj_818 (.BLUT(n2531[27]), .ALUT(n9668), .C0(n29504), .Z(n10_adj_9261));
    LUT4 i1_2_lut_3_lut_4_lut_adj_819 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(keymem_sboxw[24]), .D(n33945), .Z(n21_adj_8257)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_819.init = 16'hf0e0;
    PFUMX i25492 (.BLUT(n1_adj_8697), .ALUT(n2_adj_8696), .C0(\muxed_round_nr[1] ), 
          .Z(n30651));
    LUT4 i1_2_lut_3_lut_4_lut_adj_820 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(keymem_sboxw[25]), .D(n33945), .Z(n21_adj_8258)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_820.init = 16'hf0e0;
    PFUMX i10_adj_821 (.BLUT(n2531[28]), .ALUT(n9670), .C0(n29504), .Z(n10_adj_9264));
    PFUMX i25493 (.BLUT(n4_adj_8695), .ALUT(n5_adj_8694), .C0(\muxed_round_nr[1] ), 
          .Z(n30652));
    PFUMX i10_adj_822 (.BLUT(n2531[29]), .ALUT(n9672), .C0(n29504), .Z(n10_adj_9268));
    PFUMX i25494 (.BLUT(n8_adj_8693), .ALUT(n9_adj_8692), .C0(\muxed_round_nr[1] ), 
          .Z(n30653));
    PFUMX i10_adj_823 (.BLUT(n2531[30]), .ALUT(n9674), .C0(n29504), .Z(n10_adj_9270));
    LUT4 round_3__I_0_Mux_116_i1_3_lut (.A(\key_mem[0] [116]), .B(\key_mem[1] [116]), 
         .C(n33952), .Z(n1_adj_8708)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(178[31:36])
    defparam round_3__I_0_Mux_116_i1_3_lut.init = 16'hcaca;
    PFUMX i25499 (.BLUT(n1_adj_8690), .ALUT(n2_adj_8689), .C0(\muxed_round_nr[1] ), 
          .Z(n30658));
    PFUMX i10_adj_824 (.BLUT(n2531[31]), .ALUT(n9676), .C0(n29504), .Z(n10_adj_9272));
    LUT4 i1_2_lut_3_lut_4_lut_adj_825 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(keymem_sboxw[26]), .D(n33945), .Z(n21_adj_8259)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_825.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_826 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(keymem_sboxw[27]), .D(n33945), .Z(n21_adj_8260)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_826.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_827 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(keymem_sboxw[28]), .D(n33945), .Z(n21_adj_8261)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_827.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_828 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(keymem_sboxw[29]), .D(n33945), .Z(n21_adj_8262)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_828.init = 16'hf0e0;
    PFUMX i25500 (.BLUT(n4_adj_8688), .ALUT(n5_adj_8687), .C0(\muxed_round_nr[1] ), 
          .Z(n30659));
    FD1P3AX key_mem_ctrl_reg_FSM_i0_i1_rep_685 (.D(n6361[2]), .SP(key_mem_ctrl_we), 
            .CK(clk_c), .Q(clk_c_enable_1936));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam key_mem_ctrl_reg_FSM_i0_i1_rep_685.GSR = "ENABLED";
    FD1P3AX key_mem_ctrl_reg_FSM_i0_i1_rep_684 (.D(n6361[2]), .SP(key_mem_ctrl_we), 
            .CK(clk_c), .Q(clk_c_enable_1886));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam key_mem_ctrl_reg_FSM_i0_i1_rep_684.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_4_lut_adj_829 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[58]), .D(n33945), .Z(n22_adj_8290)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_829.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_830 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[59]), .D(n33945), .Z(n22_adj_8291)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_830.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_831 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[60]), .D(n33945), .Z(n22_adj_8292)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_831.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_832 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[61]), .D(n33945), .Z(n22_adj_8293)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_832.init = 16'hf0e0;
    FD1P3AX key_mem_ctrl_reg_FSM_i0_i1_rep_683 (.D(n6361[2]), .SP(key_mem_ctrl_we), 
            .CK(clk_c), .Q(clk_c_enable_1836));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam key_mem_ctrl_reg_FSM_i0_i1_rep_683.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_4_lut_adj_833 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[62]), .D(n33945), .Z(n22_adj_8294)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_833.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_834 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[63]), .D(n33945), .Z(n22_adj_8295)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_834.init = 16'hf0e0;
    FD1P3AX key_mem_ctrl_reg_FSM_i0_i1_rep_682 (.D(n6361[2]), .SP(key_mem_ctrl_we), 
            .CK(clk_c), .Q(clk_c_enable_1786));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam key_mem_ctrl_reg_FSM_i0_i1_rep_682.GSR = "ENABLED";
    LUT4 i14942_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[64]), .D(n33945), .Z(n8680[64])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14942_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i14943_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[65]), .D(n33945), .Z(n8680[65])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14943_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i14944_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[66]), .D(n33945), .Z(n8680[66])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14944_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i14945_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[67]), .D(n33945), .Z(n8680[67])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14945_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i14946_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[68]), .D(n33945), .Z(n8680[68])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14946_2_lut_3_lut_4_lut.init = 16'hf0e0;
    FD1P3AX key_mem_ctrl_reg_FSM_i0_i1_rep_681 (.D(n6361[2]), .SP(key_mem_ctrl_we), 
            .CK(clk_c), .Q(clk_c_enable_1736));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam key_mem_ctrl_reg_FSM_i0_i1_rep_681.GSR = "ENABLED";
    LUT4 i14947_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[69]), .D(n33945), .Z(n8680[69])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14947_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i14948_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[70]), .D(n33945), .Z(n8680[70])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14948_2_lut_3_lut_4_lut.init = 16'hf0e0;
    PFUMX i25501 (.BLUT(n8_adj_8686), .ALUT(n9_adj_8685), .C0(\muxed_round_nr[1] ), 
          .Z(n30660));
    LUT4 i14949_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[71]), .D(n33945), .Z(n8680[71])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14949_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i14950_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[72]), .D(n33945), .Z(n8680[72])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14950_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i14951_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[73]), .D(n33945), .Z(n8680[73])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14951_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i14952_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[74]), .D(n33945), .Z(n8680[74])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14952_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i14953_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[75]), .D(n33945), .Z(n8680[75])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14953_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i14954_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[76]), .D(n33945), .Z(n8680[76])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14954_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i14955_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[77]), .D(n33945), .Z(n8680[77])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14955_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i14956_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[78]), .D(n33945), .Z(n8680[78])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14956_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i14957_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[79]), .D(n33945), .Z(n8680[79])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14957_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i14958_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[80]), .D(n33945), .Z(n8680[80])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14958_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i14961_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[83]), .D(n33945), .Z(n8680[83])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14961_2_lut_3_lut_4_lut.init = 16'hf0e0;
    FD1P3AX key_mem_ctrl_reg_FSM_i0_i1_rep_680 (.D(n6361[2]), .SP(key_mem_ctrl_we), 
            .CK(clk_c), .Q(clk_c_enable_1686));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam key_mem_ctrl_reg_FSM_i0_i1_rep_680.GSR = "ENABLED";
    PFUMX i25506 (.BLUT(n1_adj_8676), .ALUT(n2_adj_8675), .C0(\muxed_round_nr[1] ), 
          .Z(n30665));
    LUT4 i14962_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[84]), .D(n33945), .Z(n8680[84])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14962_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i14965_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[87]), .D(n33945), .Z(n8680[87])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14965_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i14966_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[88]), .D(n33945), .Z(n8680[88])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14966_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i14970_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[92]), .D(n33945), .Z(n8680[92])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14970_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i14971_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[93]), .D(n33945), .Z(n8680[93])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14971_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i14973_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[95]), .D(n33945), .Z(n8680[95])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14973_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i14975_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[97]), .D(n33945), .Z(n8680[97])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14975_2_lut_3_lut_4_lut.init = 16'hf0e0;
    FD1P3AX key_mem_ctrl_reg_FSM_i0_i1_rep_679 (.D(n6361[2]), .SP(key_mem_ctrl_we), 
            .CK(clk_c), .Q(clk_c_enable_1636));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam key_mem_ctrl_reg_FSM_i0_i1_rep_679.GSR = "ENABLED";
    LUT4 i14977_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[99]), .D(n33945), .Z(n8680[99])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14977_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i14978_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[100]), .D(n33945), .Z(n8680[100])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14978_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i14980_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[102]), .D(n33945), .Z(n8680[102])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14980_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i14982_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[104]), .D(n33945), .Z(n8680[104])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14982_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i14985_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[107]), .D(n33945), .Z(n8680[107])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14985_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i14987_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[109]), .D(n33945), .Z(n8680[109])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14987_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i14989_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[111]), .D(n33945), .Z(n8680[111])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14989_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i14991_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[113]), .D(n33945), .Z(n8680[113])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14991_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i14993_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[115]), .D(n33945), .Z(n8680[115])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14993_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i14994_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[116]), .D(n33945), .Z(n8680[116])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14994_2_lut_3_lut_4_lut.init = 16'hf0e0;
    PFUMX i25507 (.BLUT(n4_adj_8649), .ALUT(n5_adj_8646), .C0(\muxed_round_nr[1] ), 
          .Z(n30666));
    LUT4 i1_2_lut_3_lut_4_lut_adj_835 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[121]), .D(n33945), .Z(n8680[121])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_835.init = 16'hf0e0;
    LUT4 i14999_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[122]), .D(n33945), .Z(n8680[122])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i14999_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i15000_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[123]), .D(n33945), .Z(n8680[123])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i15000_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i15002_2_lut_3_lut_4_lut (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[125]), .D(n33945), .Z(n8680[125])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i15002_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_836 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[126]), .D(n33945), .Z(n8680[126])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_836.init = 16'hf0e0;
    FD1P3AX key_mem_ctrl_reg_FSM_i0_i1_rep_678 (.D(n6361[2]), .SP(key_mem_ctrl_we), 
            .CK(clk_c), .Q(clk_c_enable_1586));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam key_mem_ctrl_reg_FSM_i0_i1_rep_678.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_4_lut_adj_837 (.A(round_ctr_reg[2]), .B(round_ctr_reg[3]), 
         .C(prev_key1_reg[127]), .D(n33945), .Z(n8680[127])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam i1_2_lut_3_lut_4_lut_adj_837.init = 16'hf0e0;
    LUT4 equal_138_i5_2_lut_rep_641 (.A(n35834), .B(round_ctr_reg[1]), .Z(n33945)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam equal_138_i5_2_lut_rep_641.init = 16'hdddd;
    LUT4 equal_121_i7_2_lut_rep_555_3_lut_4_lut (.A(n35834), .B(round_ctr_reg[1]), 
         .C(round_ctr_reg[3]), .D(round_ctr_reg[2]), .Z(n33859)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(157[13:35])
    defparam equal_121_i7_2_lut_rep_555_3_lut_4_lut.init = 16'hfffd;
    FD1P3AX key_mem_ctrl_reg_FSM_i0_i1_rep_677 (.D(n6361[2]), .SP(key_mem_ctrl_we), 
            .CK(clk_c), .Q(clk_c_enable_1536));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam key_mem_ctrl_reg_FSM_i0_i1_rep_677.GSR = "ENABLED";
    FD1P3AX key_mem_ctrl_reg_FSM_i0_i1_rep_676 (.D(n6361[2]), .SP(key_mem_ctrl_we), 
            .CK(clk_c), .Q(clk_c_enable_1486));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam key_mem_ctrl_reg_FSM_i0_i1_rep_676.GSR = "ENABLED";
    PFUMX i25508 (.BLUT(n8_adj_8641), .ALUT(n9_adj_8636), .C0(\muxed_round_nr[1] ), 
          .Z(n30667));
    FD1P3AX key_mem_ctrl_reg_FSM_i0_i1_rep_675 (.D(n6361[2]), .SP(key_mem_ctrl_we), 
            .CK(clk_c), .Q(clk_c_enable_1436));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam key_mem_ctrl_reg_FSM_i0_i1_rep_675.GSR = "ENABLED";
    PFUMX i25513 (.BLUT(n1_adj_8616), .ALUT(n2_adj_8611), .C0(\muxed_round_nr[1] ), 
          .Z(n30672));
    PFUMX i25514 (.BLUT(n4_adj_8604), .ALUT(n5_adj_8603), .C0(\muxed_round_nr[1] ), 
          .Z(n30673));
    FD1P3AX key_mem_ctrl_reg_FSM_i0_i1_rep_674 (.D(n6361[2]), .SP(key_mem_ctrl_we), 
            .CK(clk_c), .Q(clk_c_enable_1386));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam key_mem_ctrl_reg_FSM_i0_i1_rep_674.GSR = "ENABLED";
    PFUMX i25515 (.BLUT(n8_adj_8601), .ALUT(n9_adj_8599), .C0(\muxed_round_nr[1] ), 
          .Z(n30674));
    FD1P3AX key_mem_ctrl_reg_FSM_i0_i1_rep_673 (.D(n6361[2]), .SP(key_mem_ctrl_we), 
            .CK(clk_c), .Q(clk_c_enable_1336));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam key_mem_ctrl_reg_FSM_i0_i1_rep_673.GSR = "ENABLED";
    FD1P3AX key_mem_ctrl_reg_FSM_i0_i1_rep_672 (.D(n6361[2]), .SP(key_mem_ctrl_we), 
            .CK(clk_c), .Q(clk_c_enable_1286));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam key_mem_ctrl_reg_FSM_i0_i1_rep_672.GSR = "ENABLED";
    FD1P3AX key_mem_ctrl_reg_FSM_i0_i1_rep_671 (.D(n6361[2]), .SP(key_mem_ctrl_we), 
            .CK(clk_c), .Q(clk_c_enable_1236));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam key_mem_ctrl_reg_FSM_i0_i1_rep_671.GSR = "ENABLED";
    FD1P3AX key_mem_ctrl_reg_FSM_i0_i1_rep_670 (.D(n6361[2]), .SP(key_mem_ctrl_we), 
            .CK(clk_c), .Q(clk_c_enable_1186));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam key_mem_ctrl_reg_FSM_i0_i1_rep_670.GSR = "ENABLED";
    PFUMX i25520 (.BLUT(n1_adj_8589), .ALUT(n2_adj_8588), .C0(\muxed_round_nr[1] ), 
          .Z(n30679));
    PFUMX i25521 (.BLUT(n4_adj_8581), .ALUT(n5_adj_8577), .C0(\muxed_round_nr[1] ), 
          .Z(n30680));
    LUT4 select_751_Select_0_i4_2_lut_rep_647 (.A(\key_mem_ctrl_new_2__N_4928[0] ), 
         .B(n6361[3]), .Z(n33951)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam select_751_Select_0_i4_2_lut_rep_647.init = 16'h8888;
    LUT4 i3041_3_lut_4_lut (.A(\key_mem_ctrl_new_2__N_4928[0] ), .B(n6361[3]), 
         .C(key_ready), .D(n6361[0]), .Z(n8478)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (C+(D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam i3041_3_lut_4_lut.init = 16'hff70;
    FD1P3AX key_mem_ctrl_reg_FSM_i0_i1_rep_669 (.D(n6361[2]), .SP(key_mem_ctrl_we), 
            .CK(clk_c), .Q(clk_c_enable_1136));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam key_mem_ctrl_reg_FSM_i0_i1_rep_669.GSR = "ENABLED";
    FD1P3AX key_mem_ctrl_reg_FSM_i0_i1_rep_668 (.D(n6361[2]), .SP(key_mem_ctrl_we), 
            .CK(clk_c), .Q(clk_c_enable_1086));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam key_mem_ctrl_reg_FSM_i0_i1_rep_668.GSR = "ENABLED";
    FD1P3AX key_mem_ctrl_reg_FSM_i0_i1_rep_667 (.D(n6361[2]), .SP(key_mem_ctrl_we), 
            .CK(clk_c), .Q(clk_c_enable_1036));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam key_mem_ctrl_reg_FSM_i0_i1_rep_667.GSR = "ENABLED";
    PFUMX i25522 (.BLUT(n8_adj_8568), .ALUT(n9_adj_8567), .C0(\muxed_round_nr[1] ), 
          .Z(n30681));
    FD1P3AX key_mem_ctrl_reg_FSM_i0_i1_rep_666 (.D(n6361[2]), .SP(key_mem_ctrl_we), 
            .CK(clk_c), .Q(clk_c_enable_986));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam key_mem_ctrl_reg_FSM_i0_i1_rep_666.GSR = "ENABLED";
    FD1P3AX key_mem_ctrl_reg_FSM_i0_i1_rep_665 (.D(n6361[2]), .SP(key_mem_ctrl_we), 
            .CK(clk_c), .Q(clk_c_enable_936));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam key_mem_ctrl_reg_FSM_i0_i1_rep_665.GSR = "ENABLED";
    PFUMX i25527 (.BLUT(n1_adj_8563), .ALUT(n2_adj_8562), .C0(\muxed_round_nr[1] ), 
          .Z(n30686));
    FD1P3AX key_mem_ctrl_reg_FSM_i0_i1_rep_664 (.D(n6361[2]), .SP(key_mem_ctrl_we), 
            .CK(clk_c), .Q(clk_c_enable_886));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam key_mem_ctrl_reg_FSM_i0_i1_rep_664.GSR = "ENABLED";
    FD1P3AX key_mem_ctrl_reg_FSM_i0_i1_rep_663 (.D(n6361[2]), .SP(key_mem_ctrl_we), 
            .CK(clk_c), .Q(clk_c_enable_836));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam key_mem_ctrl_reg_FSM_i0_i1_rep_663.GSR = "ENABLED";
    LUT4 i2_4_lut_adj_838 (.A(n28850), .B(n33860), .C(\key_mem_ctrl.num_rounds[2] ), 
         .D(n33859), .Z(clk_c_enable_132)) /* synthesis lut_function=(A (B (C (D))+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam i2_4_lut_adj_838.init = 16'ha020;
    FD1P3AX key_mem_ctrl_reg_FSM_i0_i1_rep_662 (.D(n6361[2]), .SP(key_mem_ctrl_we), 
            .CK(clk_c), .Q(clk_c_enable_786));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam key_mem_ctrl_reg_FSM_i0_i1_rep_662.GSR = "ENABLED";
    PFUMX i25528 (.BLUT(n4_adj_8560), .ALUT(n5_adj_8555), .C0(\muxed_round_nr[1] ), 
          .Z(n30687));
    PFUMX i25529 (.BLUT(n8_adj_8550), .ALUT(n9_adj_8549), .C0(\muxed_round_nr[1] ), 
          .Z(n30688));
    PFUMX i25534 (.BLUT(n1_adj_8545), .ALUT(n2_adj_8542), .C0(\muxed_round_nr[1] ), 
          .Z(n30693));
    FD1P3AX key_mem_ctrl_reg_FSM_i0_i1_rep_661 (.D(n6361[2]), .SP(key_mem_ctrl_we), 
            .CK(clk_c), .Q(clk_c_enable_736));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam key_mem_ctrl_reg_FSM_i0_i1_rep_661.GSR = "ENABLED";
    PFUMX i25535 (.BLUT(n4_adj_8536), .ALUT(n5_adj_8535), .C0(\muxed_round_nr[1] ), 
          .Z(n30694));
    FD1P3AX key_mem_ctrl_reg_FSM_i0_i1_rep_660 (.D(n6361[2]), .SP(key_mem_ctrl_we), 
            .CK(clk_c), .Q(clk_c_enable_686));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam key_mem_ctrl_reg_FSM_i0_i1_rep_660.GSR = "ENABLED";
    PFUMX i25536 (.BLUT(n8_adj_8508), .ALUT(n9_adj_8502), .C0(\muxed_round_nr[1] ), 
          .Z(n30695));
    FD1P3AX key_mem_ctrl_reg_FSM_i0_i1_rep_659 (.D(n6361[2]), .SP(key_mem_ctrl_we), 
            .CK(clk_c), .Q(clk_c_enable_636));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam key_mem_ctrl_reg_FSM_i0_i1_rep_659.GSR = "ENABLED";
    FD1P3AX key_mem_ctrl_reg_FSM_i0_i1_rep_658 (.D(n6361[2]), .SP(key_mem_ctrl_we), 
            .CK(clk_c), .Q(clk_c_enable_586));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam key_mem_ctrl_reg_FSM_i0_i1_rep_658.GSR = "ENABLED";
    FD1P3AX key_mem_ctrl_reg_FSM_i0_i1_rep_657 (.D(n6361[2]), .SP(key_mem_ctrl_we), 
            .CK(clk_c), .Q(clk_c_enable_536));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam key_mem_ctrl_reg_FSM_i0_i1_rep_657.GSR = "ENABLED";
    PFUMX i25541 (.BLUT(n1_adj_8476), .ALUT(n2_adj_8473), .C0(\muxed_round_nr[1] ), 
          .Z(n30700));
    FD1P3AX key_mem_ctrl_reg_FSM_i0_i1_rep_656 (.D(n6361[2]), .SP(key_mem_ctrl_we), 
            .CK(clk_c), .Q(clk_c_enable_486));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam key_mem_ctrl_reg_FSM_i0_i1_rep_656.GSR = "ENABLED";
    FD1P3AX key_mem_ctrl_reg_FSM_i0_i1_rep_655 (.D(n6361[2]), .SP(key_mem_ctrl_we), 
            .CK(clk_c), .Q(clk_c_enable_436));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam key_mem_ctrl_reg_FSM_i0_i1_rep_655.GSR = "ENABLED";
    PFUMX i25542 (.BLUT(n4_adj_8472), .ALUT(n5_adj_8471), .C0(\muxed_round_nr[1] ), 
          .Z(n30701));
    FD1P3AX key_mem_ctrl_reg_FSM_i0_i1_rep_654 (.D(n6361[2]), .SP(key_mem_ctrl_we), 
            .CK(clk_c), .Q(n35839));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam key_mem_ctrl_reg_FSM_i0_i1_rep_654.GSR = "ENABLED";
    PFUMX i25543 (.BLUT(n8_adj_8467), .ALUT(n9_adj_8461), .C0(\muxed_round_nr[1] ), 
          .Z(n30702));
    LUT4 i15040_2_lut_4_lut (.A(\key_reg[4] [5]), .B(n4_adj_8336), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[101])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15040_2_lut_4_lut.init = 16'hca00;
    LUT4 i15039_2_lut_4_lut (.A(\key_reg[4] [4]), .B(n4_adj_8335), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[100])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15039_2_lut_4_lut.init = 16'hca00;
    LUT4 i15038_2_lut_4_lut (.A(\key_reg[4] [3]), .B(n4_adj_8333), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[99])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15038_2_lut_4_lut.init = 16'hca00;
    PFUMX i25548 (.BLUT(n1_adj_8383), .ALUT(n2_adj_8365), .C0(\muxed_round_nr[1] ), 
          .Z(n30707));
    LUT4 i15037_2_lut_4_lut (.A(\key_reg[4] [2]), .B(n4_adj_8332), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[98])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15037_2_lut_4_lut.init = 16'hca00;
    LUT4 i15036_2_lut_4_lut (.A(\key_reg[4] [1]), .B(n8929), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[97])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15036_2_lut_4_lut.init = 16'hca00;
    LUT4 i15035_2_lut_4_lut (.A(\key_reg[4] [0]), .B(n8487), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[96])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15035_2_lut_4_lut.init = 16'hca00;
    LUT4 i5_2_lut_rep_255_3_lut (.A(prev_key1_reg[95]), .B(n33716), .C(prev_key1_reg[63]), 
         .Z(n33559)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i5_2_lut_rep_255_3_lut.init = 16'h9696;
    LUT4 i3288_3_lut_4_lut (.A(prev_key1_reg[95]), .B(n33716), .C(n35835), 
         .D(n33510), .Z(n8773)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i3288_3_lut_4_lut.init = 16'hf606;
    LUT4 i6_2_lut_3_lut_4_lut (.A(prev_key1_reg[95]), .B(n33716), .C(keymem_sboxw[31]), 
         .D(prev_key1_reg[63]), .Z(n17217)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i6_2_lut_3_lut_4_lut.init = 16'h6996;
    PFUMX i25549 (.BLUT(n4_adj_8359), .ALUT(n5_adj_8356), .C0(\muxed_round_nr[1] ), 
          .Z(n30708));
    LUT4 mux_51_i96_3_lut_4_lut (.A(prev_key1_reg[95]), .B(n33716), .C(n33860), 
         .D(\key_reg[1] [31]), .Z(key_mem_new_127__N_7264[95])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam mux_51_i96_3_lut_4_lut.init = 16'h6f60;
    LUT4 i5_2_lut_rep_256_3_lut (.A(prev_key1_reg[94]), .B(n33717), .C(prev_key1_reg[62]), 
         .Z(n33560)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i5_2_lut_rep_256_3_lut.init = 16'h9696;
    LUT4 mux_51_i95_3_lut_4_lut (.A(prev_key1_reg[94]), .B(n33717), .C(n33860), 
         .D(\key_reg[1] [30]), .Z(key_mem_new_127__N_7264[94])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam mux_51_i95_3_lut_4_lut.init = 16'h6f60;
    LUT4 i6_2_lut_3_lut_4_lut_adj_839 (.A(prev_key1_reg[94]), .B(n33717), 
         .C(keymem_sboxw[30]), .D(prev_key1_reg[62]), .Z(n17157)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i6_2_lut_3_lut_4_lut_adj_839.init = 16'h6996;
    LUT4 i3286_3_lut_4_lut (.A(prev_key1_reg[94]), .B(n33717), .C(n35835), 
         .D(n33511), .Z(n8771)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i3286_3_lut_4_lut.init = 16'hf606;
    PFUMX i25550 (.BLUT(n8_adj_8350), .ALUT(n9_adj_8348), .C0(\muxed_round_nr[1] ), 
          .Z(n30709));
    LUT4 i5_2_lut_rep_259_4_lut (.A(n33718), .B(prev_key1_reg[93]), .C(prev_key1_reg[125]), 
         .D(prev_key1_reg[61]), .Z(n33563)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i5_2_lut_rep_259_4_lut.init = 16'h6996;
    LUT4 i5_2_lut_rep_260_4_lut (.A(n33719), .B(prev_key1_reg[92]), .C(prev_key1_reg[124]), 
         .D(prev_key1_reg[60]), .Z(n33564)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i5_2_lut_rep_260_4_lut.init = 16'h6996;
    LUT4 i5_2_lut_rep_262_4_lut (.A(n33720), .B(prev_key1_reg[91]), .C(prev_key1_reg[123]), 
         .D(prev_key1_reg[59]), .Z(n33566)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i5_2_lut_rep_262_4_lut.init = 16'h6996;
    PFUMX i25555 (.BLUT(n1_adj_8319), .ALUT(n2_adj_8318), .C0(\muxed_round_nr[1] ), 
          .Z(n30714));
    LUT4 i5_2_lut_rep_265_4_lut (.A(n33721), .B(prev_key1_reg[90]), .C(prev_key1_reg[122]), 
         .D(prev_key1_reg[58]), .Z(n33569)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i5_2_lut_rep_265_4_lut.init = 16'h6996;
    LUT4 i6_2_lut_3_lut_4_lut_adj_840 (.A(prev_key1_reg[89]), .B(n33722), 
         .C(keymem_sboxw[25]), .D(prev_key1_reg[57]), .Z(n16857)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i6_2_lut_3_lut_4_lut_adj_840.init = 16'h6996;
    PFUMX i25556 (.BLUT(n4_adj_8317), .ALUT(n5_adj_8316), .C0(\muxed_round_nr[1] ), 
          .Z(n30715));
    LUT4 i15025_2_lut_4_lut (.A(\key_reg[5] [22]), .B(n33623), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[86])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15025_2_lut_4_lut.init = 16'hca00;
    LUT4 i1_4_lut_adj_841 (.A(n6361[0]), .B(n6361[3]), .C(n2952), .D(\key_mem_ctrl_new_2__N_4928[0] ), 
         .Z(n28834)) /* synthesis lut_function=(A+(B (C+!(D))+!B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam i1_4_lut_adj_841.init = 16'hfafe;
    LUT4 i299_2_lut (.A(n7), .B(n35839), .Z(n2952)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(382[7] 423[14])
    defparam i299_2_lut.init = 16'h8888;
    PFUMX i25557 (.BLUT(n8_adj_8315), .ALUT(n9_adj_8308), .C0(\muxed_round_nr[1] ), 
          .Z(n30716));
    LUT4 i15024_2_lut_4_lut (.A(\key_reg[5] [21]), .B(n33625), .C(n33859), 
         .D(n33860), .Z(prev_key1_new_127__N_7520[85])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(272[19] 295[22])
    defparam i15024_2_lut_4_lut.init = 16'hca00;
    LUT4 i27845_2_lut (.A(block_w3_we_N_1490), .B(block_w2_we_N_1489), .Z(n29504)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(181[17:28])
    defparam i27845_2_lut.init = 16'heeee;
    PFUMX i25562 (.BLUT(n1_adj_8234), .ALUT(n2_adj_8233), .C0(\muxed_round_nr[1] ), 
          .Z(n30721));
    LUT4 i3276_3_lut_4_lut (.A(prev_key1_reg[89]), .B(n33722), .C(n35835), 
         .D(n33516), .Z(n8761)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i3276_3_lut_4_lut.init = 16'hf606;
    PFUMX i25563 (.BLUT(n4_adj_8232), .ALUT(n5_adj_8231), .C0(\muxed_round_nr[1] ), 
          .Z(n30722));
    LUT4 i5_2_lut_rep_266_3_lut (.A(prev_key1_reg[89]), .B(n33722), .C(prev_key1_reg[57]), 
         .Z(n33570)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i5_2_lut_rep_266_3_lut.init = 16'h9696;
    LUT4 mux_51_i90_3_lut_4_lut (.A(prev_key1_reg[89]), .B(n33722), .C(n33860), 
         .D(\key_reg[1] [25]), .Z(key_mem_new_127__N_7264[89])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam mux_51_i90_3_lut_4_lut.init = 16'h6f60;
    LUT4 i5_2_lut_rep_268_4_lut (.A(n33723), .B(prev_key1_reg[88]), .C(prev_key1_reg[120]), 
         .D(prev_key1_reg[56]), .Z(n33572)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(245[26:39])
    defparam i5_2_lut_rep_268_4_lut.init = 16'h6996;
    PFUMX i25564 (.BLUT(n8_adj_8230), .ALUT(n9_adj_8229), .C0(\muxed_round_nr[1] ), 
          .Z(n30723));
    LUT4 i6_2_lut_3_lut_adj_842 (.A(prev_key1_reg[55]), .B(n33724), .C(keymem_sboxw[23]), 
         .Z(n16737)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;
    defparam i6_2_lut_3_lut_adj_842.init = 16'h9696;
    LUT4 i2_2_lut_rep_317 (.A(prev_key0_reg[87]), .B(n4_adj_8421), .Z(n33621)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(281[23] 287[26])
    defparam i2_2_lut_rep_317.init = 16'h6666;
    PFUMX i25569 (.BLUT(n1_adj_9288), .ALUT(n2_adj_9287), .C0(\muxed_round_nr[1] ), 
          .Z(n30728));
    PFUMX i25570 (.BLUT(n4_adj_9286), .ALUT(n5_adj_9285), .C0(\muxed_round_nr[1] ), 
          .Z(n30729));
    PFUMX i25571 (.BLUT(n8_adj_9284), .ALUT(n9_adj_9283), .C0(\muxed_round_nr[1] ), 
          .Z(n30730));
    PFUMX i25576 (.BLUT(n1_adj_9281), .ALUT(n2_adj_9280), .C0(\muxed_round_nr[1] ), 
          .Z(n30735));
    PFUMX i25577 (.BLUT(n4_adj_9279), .ALUT(n5_adj_9278), .C0(\muxed_round_nr[1] ), 
          .Z(n30736));
    PFUMX i25578 (.BLUT(n8_adj_9277), .ALUT(n9_adj_9276), .C0(\muxed_round_nr[1] ), 
          .Z(n30737));
    PFUMX i25583 (.BLUT(n1_adj_9274), .ALUT(n2_adj_9273), .C0(\muxed_round_nr[1] ), 
          .Z(n30742));
    PFUMX i25584 (.BLUT(n4_adj_9271), .ALUT(n5_adj_9269), .C0(\muxed_round_nr[1] ), 
          .Z(n30743));
    PFUMX i25585 (.BLUT(n8_adj_9267), .ALUT(n9_adj_9266), .C0(\muxed_round_nr[1] ), 
          .Z(n30744));
    PFUMX i25590 (.BLUT(n1_adj_9263), .ALUT(n2_adj_9262), .C0(\muxed_round_nr[1] ), 
          .Z(n30749));
    PFUMX i25591 (.BLUT(n4_adj_9259), .ALUT(n5_adj_9257), .C0(\muxed_round_nr[1] ), 
          .Z(n30750));
    PFUMX i25592 (.BLUT(n8_adj_9255), .ALUT(n9_adj_9254), .C0(\muxed_round_nr[1] ), 
          .Z(n30751));
    PFUMX i25597 (.BLUT(n1_adj_9219), .ALUT(n2_adj_9218), .C0(\muxed_round_nr[1] ), 
          .Z(n30756));
    PFUMX i25598 (.BLUT(n4_adj_9217), .ALUT(n5_c), .C0(\muxed_round_nr[1] ), 
          .Z(n30757));
    
endmodule
//
// Verilog Description of module aes_encipher_block
//

module aes_encipher_block (n6347, clk_c, \new_sboxw[19] , n33846, \new_sboxw[20] , 
            enc_ready, n6428, \new_sboxw[21] , \round_key_gen.trw[1] , 
            round_key, \block_reg[0][5] , \round_key_gen.trw[13] , \block_reg[0][4] , 
            \round_key_gen.trw[12] , \block_reg[0][0] , \enc_new_block[56] , 
            \enc_new_block[24] , n6364, n9662, \enc_new_block[120] , 
            \enc_new_block[88] , n2531, \enc_new_block[40] , \round_key_gen.trw[8] , 
            \block_reg[1][31] , \round_key_gen.trw[3] , \enc_new_block[55] , 
            \enc_new_block[23] , n9660, \enc_new_block[119] , \enc_new_block[87] , 
            \round_logic.mixcolumns_block_71__N_1149[0] , \round_key_gen.trw[7] , 
            \round_key_gen.trw[4] , \enc_new_block[54] , \enc_new_block[22] , 
            n9658, \block_reg[1][30] , \enc_new_block[118] , \enc_new_block[86] , 
            \round_key_gen.trw[6] , \enc_new_block[53] , \enc_new_block[21] , 
            n9656, \enc_new_block[117] , \enc_new_block[85] , \round_key_gen.trw[9] , 
            \round_key_gen.trw[10] , \enc_new_block[52] , \enc_new_block[20] , 
            n9654, \block_reg[1][29] , \enc_new_block[116] , \enc_new_block[84] , 
            \enc_new_block[51] , \enc_new_block[19] , n9652, \round_key_gen.trw[5] , 
            \enc_new_block[115] , \enc_new_block[83] , \round_key_gen.trw[11] , 
            \enc_new_block[50] , \enc_new_block[18] , n9650, \enc_new_block[58] , 
            \round_key_gen.trw[14] , \round_key_gen.trw[17] , \block_reg[1][26] , 
            \enc_new_block[114] , \enc_new_block[82] , \round_key_gen.trw[19] , 
            \enc_new_block[49] , \enc_new_block[17] , n9648, \enc_new_block[67] , 
            \enc_new_block[113] , \enc_new_block[81] , \round_key_gen.trw[20] , 
            \enc_new_block[48] , \enc_new_block[16] , n9646, \enc_new_block[112] , 
            \enc_new_block[80] , \round_logic.mixcolumns_block_111__N_1285[0] , 
            \round_logic.mixcolumns_block_79__N_1341[0] , n9644, \round_logic.mixcolumns_block_47__N_1397[0] , 
            \round_logic.mixcolumns_block_15__N_1453[0] , \round_logic.mixcolumns_block_111__N_1285[7] , 
            \round_logic.mixcolumns_block_79__N_1341[7] , n9642, \round_logic.mixcolumns_block_47__N_1397[7] , 
            \round_logic.mixcolumns_block_15__N_1453[7] , \new_sboxw[17] , 
            \round_logic.mixcolumns_block_111__N_1285[6] , \round_logic.mixcolumns_block_79__N_1341[6] , 
            n9640, \new_sboxw[18] , \round_key_gen.trw[15] , \new_sboxw[22] , 
            \new_sboxw[23] , \enc_new_block[57] , \round_logic.mixcolumns_block_39__N_1197[2] , 
            \round_logic.mixcolumns_block_47__N_1397[6] , \round_logic.mixcolumns_block_15__N_1453[6] , 
            \round_logic.mixcolumns_block_111__N_1285[5] , \round_logic.mixcolumns_block_79__N_1341[5] , 
            n9638, \enc_new_block[32] , \round_logic.mixcolumns_block_7__N_1245[7] , 
            \round_logic.mixcolumns_block_47__N_1397[5] , \round_logic.mixcolumns_block_15__N_1453[5] , 
            \enc_new_block[43] , \enc_new_block[11] , n9636, \enc_new_block[107] , 
            \enc_new_block[75] , \enc_new_block[72] , \round_logic.mixcolumns_block_15__N_1453[2] , 
            \enc_new_block[42] , \enc_new_block[10] , n9634, \enc_new_block[106] , 
            \enc_new_block[74] , \round_logic.mixcolumns_block_111__N_1285[2] , 
            \round_logic.mixcolumns_block_79__N_1341[2] , n9632, \round_logic.mixcolumns_block_47__N_1397[2] , 
            \round_key_gen.trw[2] , \enc_new_block[26] , \enc_new_block[8] , 
            n9630, \enc_new_block[104] , \enc_new_block[29] , \round_logic.mixcolumns_block_7__N_1245[0] , 
            \round_logic.mixcolumns_block_103__N_1101[0] , n9628, \enc_new_block[31] , 
            \enc_new_block[64] , \round_logic.mixcolumns_block_39__N_1197[0] , 
            \round_logic.mixcolumns_block_39__N_1197[7] , \round_logic.mixcolumns_block_103__N_1101[7] , 
            n9626, \round_logic.mixcolumns_block_71__N_1149[7] , \round_logic.mixcolumns_block_7__N_1245[6] , 
            \round_logic.mixcolumns_block_103__N_1101[6] , n9624, \round_logic.mixcolumns_block_71__N_1149[6] , 
            \round_logic.mixcolumns_block_39__N_1197[6] , \round_logic.mixcolumns_block_7__N_1245[5] , 
            \round_logic.mixcolumns_block_103__N_1101[5] , n9622, \round_logic.mixcolumns_block_71__N_1149[5] , 
            \round_logic.mixcolumns_block_39__N_1197[5] , \enc_new_block[35] , 
            \enc_new_block[3] , n9620, \enc_new_block[99] , \enc_new_block[34] , 
            \enc_new_block[2] , n9618, \enc_new_block[98] , \enc_new_block[66] , 
            \round_logic.mixcolumns_block_7__N_1245[2] , \round_logic.mixcolumns_block_103__N_1101[2] , 
            n9616, \enc_new_block[63] , \round_logic.mixcolumns_block_71__N_1149[2] , 
            \enc_new_block[0] , n8532, \enc_new_block[96] , \enc_new_block[90] , 
            \enc_new_block[93] , \enc_new_block[94] , \enc_new_block[95] , 
            \enc_new_block[122] , \enc_new_block[27] , \enc_new_block[28] , 
            \enc_new_block[30] , \block_reg[0][31] , \enc_new_block[59] , 
            \enc_new_block[60] , \enc_new_block[61] , \enc_new_block[62] , 
            \block_reg[0][30] , \block_reg[0][28] , \block_reg[0][26] , 
            \enc_new_block[89] , \enc_new_block[91] , \enc_new_block[92] , 
            block_w2_we_N_1489, \block_reg[0][24] , \round_key_gen.trw[0] , 
            \block_reg[0][21] , \enc_new_block[125] , \block_reg[0][16] , 
            \new_sboxw[16] , \block_reg[0][15] , \enc_new_block[127] , 
            \round_key_gen.trw[23] , \block_reg[0][14] , \round_key_gen.trw[22] , 
            \block_reg[0][13] , \round_key_gen.trw[21] , \block_reg[0][10] , 
            \round_key_gen.trw[18] , \block_reg[0][8] , \round_key_gen.trw[16] , 
            \block_reg[0][7] , n9676, n9674, \enc_new_block[126] , n9672, 
            n9670, \enc_new_block[124] , n9668, \enc_new_block[123] , 
            n9666, \enc_new_block[25] , n9664, \enc_new_block[121] , 
            \block_new_127__N_1645[125] , \block_new_127__N_1645[123] , 
            \block_new_127__N_1645[121] , \block_new_127__N_1645[119] , 
            \block_reg[1][24] , \block_new_127__N_1645[118] , \block_new_127__N_1645[116] , 
            \block_new_127__N_1645[115] , \block_new_127__N_1645[114] , 
            \block_new_127__N_1645[113] , \block_new_127__N_1645[108] , 
            \block_reg[1][16] , \block_reg[1][15] , n33848, \block_reg[1][14] , 
            \block_reg[1][13] , \block_new_127__N_1645[107] , \block_new_127__N_1645[105] , 
            \block_new_127__N_1645[102] , \block_reg[1][10] , \block_new_127__N_1645[99] , 
            \block_new_127__N_1645[98] , \block_new_127__N_1645[97] , \block_reg[1][8] , 
            \block_reg[2][3] , enc_round_nr, \block_new_127__N_1645[92] , 
            \block_new_127__N_1645[91] , \block_new_127__N_1645[89] , \block_new_127__N_1645[87] , 
            \block_new_127__N_1645[86] , \block_new_127__N_1645[85] , \block_new_127__N_1645[84] , 
            \block_reg[1][2] , \block_new_127__N_1645[83] , \block_new_127__N_1645[82] , 
            \block_new_127__N_1645[81] , \block_new_127__N_1645[76] , \block_reg[2][31] , 
            \block_new_127__N_1645[75] , \block_new_127__N_1645[73] , \block_new_127__N_1645[71] , 
            \block_new_127__N_1645[70] , \block_reg[2][26] , n33913, n28773, 
            \block_reg[2][24] , \block_reg[2][23] , \block_new_127__N_1645[69] , 
            \block_reg[2][22] , \block_reg[2][21] , \block_reg[2][20] , 
            \block_reg[2][16] , \block_reg[2][15] , \block_reg[2][14] , 
            \block_new_127__N_1645[68] , \block_new_127__N_1645[67] , \block_reg[2][13] , 
            \block_new_127__N_1645[65] , \block_reg[2][10] , \block_new_127__N_1645[64] , 
            \block_reg[2][8] , \block_reg[2][6] , n5, round_ctr_we, 
            n33915, \block_new_127__N_1645[62] , \block_new_127__N_1645[61] , 
            \key_mem_ctrl.num_rounds[2] , n4, \block_new_127__N_1645[12] , 
            \block_new_127__N_1645[60] , \block_new_127__N_1645[10] , \block_new_127__N_1645[7] , 
            \block_new_127__N_1645[59] , \block_new_127__N_1645[5] , \block_new_127__N_1645[4] , 
            \block_new_127__N_1645[57] , \block_reg[2][0] , \block_reg[3][31] , 
            \block_reg[3][29] , \block_new_127__N_1645[3] , \block_new_127__N_1645[2] , 
            \block_reg[3][26] , \block_new_127__N_1645[1] , \block_reg[3][24] , 
            \block_reg[3][23] , \block_new_127__N_1645[51] , \block_reg[3][22] , 
            \block_new_127__N_1645[50] , \block_new_127__N_1645[49] , \block_reg[3][18] , 
            \block_new_127__N_1645[44] , \block_new_127__N_1645[43] , \block_new_127__N_1645[41] , 
            \block_reg[3][16] , \block_reg[3][15] , \block_new_127__N_1645[39] , 
            \block_new_127__N_1645[37] , \block_new_127__N_1645[36] , \block_new_127__N_1645[34] , 
            \block_reg[3][13] , \block_new_127__N_1645[33] , \block_new_127__N_1645[30] , 
            \block_reg[3][11] , \block_new_127__N_1645[28] , \block_new_127__N_1645[27] , 
            \block_reg[3][9] , \block_new_127__N_1645[25] , \block_reg[3][8] , 
            \block_reg[3][6] , \block_new_127__N_1645[21] , \block_new_127__N_1645[20] , 
            \block_new_127__N_1645[19] , \block_new_127__N_1645[17] , \block_new_127__N_1645[14] , 
            \block_reg[3][0] ) /* synthesis syn_module_defined=1 */ ;
    output [3:0]n6347;
    input clk_c;
    input \new_sboxw[19] ;
    input n33846;
    input \new_sboxw[20] ;
    output enc_ready;
    input n6428;
    input \new_sboxw[21] ;
    input \round_key_gen.trw[1] ;
    input [127:0]round_key;
    input \block_reg[0][5] ;
    input \round_key_gen.trw[13] ;
    input \block_reg[0][4] ;
    input \round_key_gen.trw[12] ;
    input \block_reg[0][0] ;
    output \enc_new_block[56] ;
    output \enc_new_block[24] ;
    output [3:0]n6364;
    output n9662;
    output \enc_new_block[120] ;
    output \enc_new_block[88] ;
    output [31:0]n2531;
    output \enc_new_block[40] ;
    input \round_key_gen.trw[8] ;
    input \block_reg[1][31] ;
    input \round_key_gen.trw[3] ;
    output \enc_new_block[55] ;
    output \enc_new_block[23] ;
    output n9660;
    output \enc_new_block[119] ;
    output \enc_new_block[87] ;
    output \round_logic.mixcolumns_block_71__N_1149[0] ;
    input \round_key_gen.trw[7] ;
    input \round_key_gen.trw[4] ;
    output \enc_new_block[54] ;
    output \enc_new_block[22] ;
    output n9658;
    input \block_reg[1][30] ;
    output \enc_new_block[118] ;
    output \enc_new_block[86] ;
    input \round_key_gen.trw[6] ;
    output \enc_new_block[53] ;
    output \enc_new_block[21] ;
    output n9656;
    output \enc_new_block[117] ;
    output \enc_new_block[85] ;
    input \round_key_gen.trw[9] ;
    input \round_key_gen.trw[10] ;
    output \enc_new_block[52] ;
    output \enc_new_block[20] ;
    output n9654;
    input \block_reg[1][29] ;
    output \enc_new_block[116] ;
    output \enc_new_block[84] ;
    output \enc_new_block[51] ;
    output \enc_new_block[19] ;
    output n9652;
    input \round_key_gen.trw[5] ;
    output \enc_new_block[115] ;
    output \enc_new_block[83] ;
    input \round_key_gen.trw[11] ;
    output \enc_new_block[50] ;
    output \enc_new_block[18] ;
    output n9650;
    output \enc_new_block[58] ;
    input \round_key_gen.trw[14] ;
    input \round_key_gen.trw[17] ;
    input \block_reg[1][26] ;
    output \enc_new_block[114] ;
    output \enc_new_block[82] ;
    input \round_key_gen.trw[19] ;
    output \enc_new_block[49] ;
    output \enc_new_block[17] ;
    output n9648;
    output \enc_new_block[67] ;
    output \enc_new_block[113] ;
    output \enc_new_block[81] ;
    input \round_key_gen.trw[20] ;
    output \enc_new_block[48] ;
    output \enc_new_block[16] ;
    output n9646;
    output \enc_new_block[112] ;
    output \enc_new_block[80] ;
    output \round_logic.mixcolumns_block_111__N_1285[0] ;
    output \round_logic.mixcolumns_block_79__N_1341[0] ;
    output n9644;
    output \round_logic.mixcolumns_block_47__N_1397[0] ;
    output \round_logic.mixcolumns_block_15__N_1453[0] ;
    output \round_logic.mixcolumns_block_111__N_1285[7] ;
    output \round_logic.mixcolumns_block_79__N_1341[7] ;
    output n9642;
    output \round_logic.mixcolumns_block_47__N_1397[7] ;
    output \round_logic.mixcolumns_block_15__N_1453[7] ;
    input \new_sboxw[17] ;
    output \round_logic.mixcolumns_block_111__N_1285[6] ;
    output \round_logic.mixcolumns_block_79__N_1341[6] ;
    output n9640;
    input \new_sboxw[18] ;
    input \round_key_gen.trw[15] ;
    input \new_sboxw[22] ;
    input \new_sboxw[23] ;
    output \enc_new_block[57] ;
    output \round_logic.mixcolumns_block_39__N_1197[2] ;
    output \round_logic.mixcolumns_block_47__N_1397[6] ;
    output \round_logic.mixcolumns_block_15__N_1453[6] ;
    output \round_logic.mixcolumns_block_111__N_1285[5] ;
    output \round_logic.mixcolumns_block_79__N_1341[5] ;
    output n9638;
    output \enc_new_block[32] ;
    output \round_logic.mixcolumns_block_7__N_1245[7] ;
    output \round_logic.mixcolumns_block_47__N_1397[5] ;
    output \round_logic.mixcolumns_block_15__N_1453[5] ;
    output \enc_new_block[43] ;
    output \enc_new_block[11] ;
    output n9636;
    output \enc_new_block[107] ;
    output \enc_new_block[75] ;
    output \enc_new_block[72] ;
    output \round_logic.mixcolumns_block_15__N_1453[2] ;
    output \enc_new_block[42] ;
    output \enc_new_block[10] ;
    output n9634;
    output \enc_new_block[106] ;
    output \enc_new_block[74] ;
    output \round_logic.mixcolumns_block_111__N_1285[2] ;
    output \round_logic.mixcolumns_block_79__N_1341[2] ;
    output n9632;
    output \round_logic.mixcolumns_block_47__N_1397[2] ;
    input \round_key_gen.trw[2] ;
    output \enc_new_block[26] ;
    output \enc_new_block[8] ;
    output n9630;
    output \enc_new_block[104] ;
    output \enc_new_block[29] ;
    output \round_logic.mixcolumns_block_7__N_1245[0] ;
    output \round_logic.mixcolumns_block_103__N_1101[0] ;
    output n9628;
    output \enc_new_block[31] ;
    output \enc_new_block[64] ;
    output \round_logic.mixcolumns_block_39__N_1197[0] ;
    output \round_logic.mixcolumns_block_39__N_1197[7] ;
    output \round_logic.mixcolumns_block_103__N_1101[7] ;
    output n9626;
    output \round_logic.mixcolumns_block_71__N_1149[7] ;
    output \round_logic.mixcolumns_block_7__N_1245[6] ;
    output \round_logic.mixcolumns_block_103__N_1101[6] ;
    output n9624;
    output \round_logic.mixcolumns_block_71__N_1149[6] ;
    output \round_logic.mixcolumns_block_39__N_1197[6] ;
    output \round_logic.mixcolumns_block_7__N_1245[5] ;
    output \round_logic.mixcolumns_block_103__N_1101[5] ;
    output n9622;
    output \round_logic.mixcolumns_block_71__N_1149[5] ;
    output \round_logic.mixcolumns_block_39__N_1197[5] ;
    output \enc_new_block[35] ;
    output \enc_new_block[3] ;
    output n9620;
    output \enc_new_block[99] ;
    output \enc_new_block[34] ;
    output \enc_new_block[2] ;
    output n9618;
    output \enc_new_block[98] ;
    output \enc_new_block[66] ;
    output \round_logic.mixcolumns_block_7__N_1245[2] ;
    output \round_logic.mixcolumns_block_103__N_1101[2] ;
    output n9616;
    output \enc_new_block[63] ;
    output \round_logic.mixcolumns_block_71__N_1149[2] ;
    output \enc_new_block[0] ;
    output n8532;
    output \enc_new_block[96] ;
    output \enc_new_block[90] ;
    output \enc_new_block[93] ;
    output \enc_new_block[94] ;
    output \enc_new_block[95] ;
    output \enc_new_block[122] ;
    output \enc_new_block[27] ;
    output \enc_new_block[28] ;
    output \enc_new_block[30] ;
    input \block_reg[0][31] ;
    output \enc_new_block[59] ;
    output \enc_new_block[60] ;
    output \enc_new_block[61] ;
    output \enc_new_block[62] ;
    input \block_reg[0][30] ;
    input \block_reg[0][28] ;
    input \block_reg[0][26] ;
    output \enc_new_block[89] ;
    output \enc_new_block[91] ;
    output \enc_new_block[92] ;
    output block_w2_we_N_1489;
    input \block_reg[0][24] ;
    input \round_key_gen.trw[0] ;
    input \block_reg[0][21] ;
    output \enc_new_block[125] ;
    input \block_reg[0][16] ;
    input \new_sboxw[16] ;
    input \block_reg[0][15] ;
    output \enc_new_block[127] ;
    input \round_key_gen.trw[23] ;
    input \block_reg[0][14] ;
    input \round_key_gen.trw[22] ;
    input \block_reg[0][13] ;
    input \round_key_gen.trw[21] ;
    input \block_reg[0][10] ;
    input \round_key_gen.trw[18] ;
    input \block_reg[0][8] ;
    input \round_key_gen.trw[16] ;
    input \block_reg[0][7] ;
    output n9676;
    output n9674;
    output \enc_new_block[126] ;
    output n9672;
    output n9670;
    output \enc_new_block[124] ;
    output n9668;
    output \enc_new_block[123] ;
    output n9666;
    output \enc_new_block[25] ;
    output n9664;
    output \enc_new_block[121] ;
    input \block_new_127__N_1645[125] ;
    input \block_new_127__N_1645[123] ;
    input \block_new_127__N_1645[121] ;
    input \block_new_127__N_1645[119] ;
    input \block_reg[1][24] ;
    input \block_new_127__N_1645[118] ;
    input \block_new_127__N_1645[116] ;
    input \block_new_127__N_1645[115] ;
    input \block_new_127__N_1645[114] ;
    input \block_new_127__N_1645[113] ;
    input \block_new_127__N_1645[108] ;
    input \block_reg[1][16] ;
    input \block_reg[1][15] ;
    output n33848;
    input \block_reg[1][14] ;
    input \block_reg[1][13] ;
    input \block_new_127__N_1645[107] ;
    input \block_new_127__N_1645[105] ;
    input \block_new_127__N_1645[102] ;
    input \block_reg[1][10] ;
    input \block_new_127__N_1645[99] ;
    input \block_new_127__N_1645[98] ;
    input \block_new_127__N_1645[97] ;
    input \block_reg[1][8] ;
    input \block_reg[2][3] ;
    output [3:0]enc_round_nr;
    input \block_new_127__N_1645[92] ;
    input \block_new_127__N_1645[91] ;
    input \block_new_127__N_1645[89] ;
    input \block_new_127__N_1645[87] ;
    input \block_new_127__N_1645[86] ;
    input \block_new_127__N_1645[85] ;
    input \block_new_127__N_1645[84] ;
    input \block_reg[1][2] ;
    input \block_new_127__N_1645[83] ;
    input \block_new_127__N_1645[82] ;
    input \block_new_127__N_1645[81] ;
    input \block_new_127__N_1645[76] ;
    input \block_reg[2][31] ;
    input \block_new_127__N_1645[75] ;
    input \block_new_127__N_1645[73] ;
    input \block_new_127__N_1645[71] ;
    input \block_new_127__N_1645[70] ;
    input \block_reg[2][26] ;
    input n33913;
    input n28773;
    input \block_reg[2][24] ;
    input \block_reg[2][23] ;
    input \block_new_127__N_1645[69] ;
    input \block_reg[2][22] ;
    input \block_reg[2][21] ;
    input \block_reg[2][20] ;
    input \block_reg[2][16] ;
    input \block_reg[2][15] ;
    input \block_reg[2][14] ;
    input \block_new_127__N_1645[68] ;
    input \block_new_127__N_1645[67] ;
    input \block_reg[2][13] ;
    input \block_new_127__N_1645[65] ;
    input \block_reg[2][10] ;
    input \block_new_127__N_1645[64] ;
    input \block_reg[2][8] ;
    input \block_reg[2][6] ;
    output n5;
    input round_ctr_we;
    output n33915;
    input \block_new_127__N_1645[62] ;
    input \block_new_127__N_1645[61] ;
    input \key_mem_ctrl.num_rounds[2] ;
    output n4;
    input \block_new_127__N_1645[12] ;
    input \block_new_127__N_1645[60] ;
    input \block_new_127__N_1645[10] ;
    input \block_new_127__N_1645[7] ;
    input \block_new_127__N_1645[59] ;
    input \block_new_127__N_1645[5] ;
    input \block_new_127__N_1645[4] ;
    input \block_new_127__N_1645[57] ;
    input \block_reg[2][0] ;
    input \block_reg[3][31] ;
    input \block_reg[3][29] ;
    input \block_new_127__N_1645[3] ;
    input \block_new_127__N_1645[2] ;
    input \block_reg[3][26] ;
    input \block_new_127__N_1645[1] ;
    input \block_reg[3][24] ;
    input \block_reg[3][23] ;
    input \block_new_127__N_1645[51] ;
    input \block_reg[3][22] ;
    input \block_new_127__N_1645[50] ;
    input \block_new_127__N_1645[49] ;
    input \block_reg[3][18] ;
    input \block_new_127__N_1645[44] ;
    input \block_new_127__N_1645[43] ;
    input \block_new_127__N_1645[41] ;
    input \block_reg[3][16] ;
    input \block_reg[3][15] ;
    input \block_new_127__N_1645[39] ;
    input \block_new_127__N_1645[37] ;
    input \block_new_127__N_1645[36] ;
    input \block_new_127__N_1645[34] ;
    input \block_reg[3][13] ;
    input \block_new_127__N_1645[33] ;
    input \block_new_127__N_1645[30] ;
    input \block_reg[3][11] ;
    input \block_new_127__N_1645[28] ;
    input \block_new_127__N_1645[27] ;
    input \block_reg[3][9] ;
    input \block_new_127__N_1645[25] ;
    input \block_reg[3][8] ;
    input \block_reg[3][6] ;
    input \block_new_127__N_1645[21] ;
    input \block_new_127__N_1645[20] ;
    input \block_new_127__N_1645[19] ;
    input \block_new_127__N_1645[17] ;
    input \block_new_127__N_1645[14] ;
    input \block_reg[3][0] ;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(41[33:36])
    
    wire enc_ctrl_we, n1, n7, n8, n2, n7_adj_8025, n8_adj_8026, 
        n2_adj_8027, n7_adj_8028, n8_adj_8029, n2_adj_8030, n9, n10, 
        n2_adj_8031, n32300, n32302, n32303, n32306, n28933, n33897, 
        n33893, n32308, n32309, n7_adj_8032, n8_adj_8033, n2_adj_8034, 
        n33847, n33845, n33036, n33038, n33039, n32321, n33054, 
        n33056, n33057, n33069, n33071, n33072, n33078, n33080, 
        n33081, n33090, n33092, n33093;
    wire [3:0]n6364_c;
    
    wire n33898, n32323, n32324, n32327, n7_adj_8035, n8_adj_8036, 
        n2_adj_8037, n33109, n33111, n33112, n33123, n33125, n33126, 
        n33132, n33134, n33135, n33889, n33890, n32329, n32330, 
        n7_adj_8038, n8_adj_8039, n2_adj_8040, n32333, n7_adj_8041, 
        n8_adj_8042, n2_adj_8043, n33887, n33888, n32335, n9_adj_8044, 
        n10_adj_8045, n2_adj_8046, n32336, n7_adj_8047, n8_adj_8048, 
        n2_adj_8049, n7_adj_8050, n8_adj_8051, n2_adj_8052, n7_adj_8053, 
        n8_adj_8054, n2_adj_8055, n32339, n7_adj_8056, n8_adj_8057, 
        n2_adj_8058, n33138, n33140, n33141, n33885, n33886, n32341, 
        n33159, n33161, n33162, n33173, n33175, n33176, n32342, 
        n7_adj_8059, n8_adj_8060, n2_adj_8061, n7_adj_8062, n8_adj_8063, 
        n2_adj_8064, n7_adj_8065, n8_adj_8066, n2_adj_8067, n33867, 
        n7_adj_8068, n8_adj_8069, n2_adj_8070, n7_adj_8071, n8_adj_8072, 
        n2_adj_8073, n32363, n33182, n33184, n33185, n33194, n33196, 
        n33197, n33206, n33208, n33209, n7_adj_8074, n8_adj_8075, 
        n2_adj_8076, n7_adj_8077, n9_adj_8078, n10_adj_8079, n2_adj_8080, 
        n33218, n33220, n33221, n33224, n33226, n33227, n33236, 
        n33238, n33239, n7_adj_8081, n8_adj_8082, n2_adj_8083, n33271, 
        n33273, n33274, n7_adj_8084, n8_adj_8085, n2_adj_8086, n7_adj_8087, 
        n8_adj_8088, n2_adj_8089, n7_adj_8090, n8_adj_8091, n2_adj_8092, 
        n9_adj_8093, n10_adj_8094, n2_adj_8095, n7_adj_8096, n8_adj_8097, 
        n2_adj_8098, n7_adj_8099, n8_adj_8100, n2_adj_8101, n7_adj_8102, 
        n8_adj_8103, n2_adj_8104, n7_adj_8105, n8_adj_8106, n2_adj_8107, 
        n7_adj_8108, n8_adj_8109, n2_adj_8110, n7_adj_8111, n8_adj_8112, 
        n2_adj_8113, n7_adj_8114, n8_adj_8115, n2_adj_8116, n33270, 
        n33269, n7_adj_8117, n8_adj_8118, n2_adj_8119, n33234, n33222, 
        n33878, n33879, n32365, n33216, n33204, n33192, n33180, 
        n33171, n33157, n33136, n7_adj_8120, n8_adj_8121, n2_adj_8122, 
        n33130, n32366, n33121, n33107, n33088, n33076, n33067, 
        n33052, n33034, n10_adj_8123, n33055, n33022, n33010, n32993, 
        n32984, n32978, n32969, n32948, n32939, n32933, n33868, 
        n8_adj_8124, n32919, n32909, n32896, n32850, n32784, n32697, 
        n32600, n32577, n32571, n32560, n32554, n32508, n32362, 
        n32338, n32332, n32326, n32320, n32305, n32299, n32290, 
        n32284, n32275, n32261, n32255, n32249, n32243, n32223, 
        n32211, n32202, n12960, n12961, block_w3_we, n12963, n12966, 
        n12967, n12969, n12970, n12972, n7_adj_8125, n8_adj_8126, 
        n2_adj_8127, n12974, n12976, n12977, n7_adj_8128, n8_adj_8129, 
        n2_adj_8130, n7_adj_8131, n8_adj_8132, n2_adj_8133, n12982, 
        n12983, n33235, n12984, n12990, n32177, n29399, n33908, 
        n32179, n32180, block_w0_we, n32325, n12992, n12993, n12994, 
        n12995, n32183, n12997, n12998, n13000, n13001, n33906, 
        n33907, n32185, n13002, n32186, n7_adj_8134, n8_adj_8135, 
        n2_adj_8136, n33223, n28939, n8_adj_8137, n32194, n2_adj_8138, 
        n33903, n33904, n32196, n13003, n7_adj_8139, n2_adj_8140, 
        n32197, n33217, n7_adj_8141, n8_adj_8142, n2_adj_8143, n7_adj_8144, 
        n8_adj_8145, n2_adj_8146, n32203, n33900, n33901, n32205, 
        n32206, n13004, block_w1_we;
    wire [127:0]n5291;
    
    wire n7_adj_8147, n8_adj_8148, n2_adj_8149, n33205, n13006, n13008, 
        n7_adj_8150, n8_adj_8151, n2_adj_8152, n13009, n13014, n13015, 
        n13016, n13017, n13018, n13019, n13020, n33193, n33869, 
        n13022, n13024, n13025, block_w2_we, n33841, n20690, n13030, 
        n13031, n13032, sword_ctr_we, n25323, n13035, n13038, n13040, 
        n33181, n13041, n13046, n32212, n9_adj_8153, n10_adj_8154, 
        n2_adj_8155, n29077, n32214, n7_adj_8156, n8_adj_8157, n2_adj_8158, 
        n32215, n33172, n13047, n13048, n7_adj_8159, n8_adj_8160, 
        n2_adj_8161, n7_adj_8162, n8_adj_8163, n2_adj_8164, n32178, 
        n32181, n32184, n32187, n32195, n32198, n7_adj_8165, n8_adj_8166, 
        n2_adj_8167, n32204, n32207, n32213, n32216, n32225, n32227, 
        n32228, n32245, n32247, n32248, n32251, n32253, n32254, 
        n7_adj_8168, n8_adj_8169, n2_adj_8170, n32257, n32259, n32260, 
        n32263, n32265, n32266, n32224, n33902, n29303, n32226, 
        n32277, n32279, n32280, n32286, n32288, n32289, n32292, 
        n32294, n32295, n32301, n32304, n32307, n32310, n32322, 
        n32328, n32331, n32334, n32337, n32340, n32343, n32364, 
        n32367, n32510, n32512, n32513, n32556, n32558, n32559, 
        n32562, n32564, n32565, n32573, n32575, n32576, n32579, 
        n32581, n32582, n32602, n32604, n32605, n32244, n33895, 
        n33896, n32246, n32250, n32252, n32256, n29037, n32258, 
        n32262, n33852, n32264, n32276, n33891, n33892, n32278, 
        n32285, n32287, n32291, n32699, n32701, n32702, n7_adj_8171, 
        n8_adj_8172, n2_adj_8173, n7_adj_8174, n8_adj_8175, n2_adj_8176, 
        n32786, n32788, n32789, n32852, n32854, n32855, n32898, 
        n32900, n32901, n32911, n32913, n32914, n32921, n32923, 
        n32924, n32935, n32937, n32938, n32293, n7_adj_8177, n8_adj_8178, 
        n2_adj_8179, n32941, n32943, n32944, n32950, n32952, n32953, 
        n32971, n32973, n32974, n32980, n32982, n32983, n7_adj_8180, 
        n8_adj_8181, n2_adj_8182, n7_adj_8183, n8_adj_8184, n2_adj_8185, 
        n32986, n32988, n32989, n32995, n32997, n32998, n7_adj_8186, 
        n8_adj_8187, n2_adj_8188, n33012, n33014, n33015, n33024, 
        n33026, n33027, n7_adj_8189, n8_adj_8190, n2_adj_8191, n7_adj_8192, 
        n8_adj_8193, n2_adj_8194, n7_adj_8195, n8_adj_8196, n2_adj_8197, 
        n33158, n33870, n13049, n13051, n13052, n13054, n13056, 
        n32182, n32193, n32176, n12934, n12935, n12936, n12937, 
        n12938, n12940, n12943, n12945, n12947, n12950, n12952, 
        n12953, n12954, n12958, n13058, n33871, n32511, n33137, 
        n33131, n33872, n33122, n33108, n33882, n29058;
    wire [127:0]n5932;
    
    wire n32509, n33089, n33077, n32555, n32557, n32561, n28866, 
        n32563, n32572, n32574, n32578, n33883, n32580, n32601, 
        n32603, n33068, n32698, n33875, n32700, n33053, n33914, 
        n2924, n33843, n32785, n33881, n33876, n33851, n32787, 
        n29071, n32851, n33862, n11620, n32853, n33880, n33894, 
        n33905, n11634, n11641, n11630, n33926, n12156, n29080, 
        n10_adj_8198, n7_adj_8199, n10_adj_8200, n7_adj_8201, n7_adj_8202, 
        n32897, n7_adj_8203, n33877, n7_adj_8204, n7_adj_8205, n7_adj_8206, 
        n9_adj_8207, n33922, n10_adj_8208, n29083, n33884, n29105, 
        n33899, n11593, n33866, n32899, n32910, n33863, n32912, 
        n20693, n32920, n33035, n29123, n32922, n32934, n28869, 
        n32936, n32940, n33855, n32942, n32949, n33854, n32951, 
        n32970, n33933, n32972, n32979, n32981, n32985, n32987, 
        n32994, n32996, n33011, n33864, n33013, n33023, n33025, 
        n2_adj_8209, n8_adj_8210, n2_adj_8211, n8_adj_8212, n2_adj_8213, 
        n8_adj_8214, n2_adj_8215, n8_adj_8216, n2_adj_8217, n8_adj_8218, 
        n2_adj_8219, n8_adj_8220, n2_adj_8221, n7_adj_8222, n8_adj_8223, 
        n2_adj_8224, n8_adj_8225, n2_adj_8226, n9_adj_8227, n2_adj_8228;
    wire [3:0]n21;
    
    wire n28860, n28861, n33929, n33225, n33924, n33865, n33934, 
        n33931, n33037, n33932, n33917, n33918, n33920, n33919, 
        n33921, n28930, n33925, n33923, n33927, n33928, n33853, 
        n33207, n33930, n33070, n33079, n33091, n33110, n33124, 
        n33133, n20687, n33139, n33160, n33174, n33183, n33195, 
        n20696, n33219, n33237, n33272;
    
    FD1P3AX enc_ctrl_reg_FSM_i0_i0 (.D(n1), .SP(enc_ctrl_we), .CK(clk_c), 
            .Q(n6347[0]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(422[7] 479[14])
    defparam enc_ctrl_reg_FSM_i0_i0.GSR = "ENABLED";
    LUT4 mux_692_Mux_19_i2_4_lut (.A(\new_sboxw[19] ), .B(n7), .C(n33846), 
         .D(n8), .Z(n2)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_19_i2_4_lut.init = 16'h3aca;
    LUT4 mux_692_Mux_20_i2_4_lut (.A(\new_sboxw[20] ), .B(n7_adj_8025), 
         .C(n33846), .D(n8_adj_8026), .Z(n2_adj_8027)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_20_i2_4_lut.init = 16'h3aca;
    FD1S3AY ready_reg_218 (.D(n6428), .CK(clk_c), .Q(enc_ready));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam ready_reg_218.GSR = "ENABLED";
    LUT4 mux_692_Mux_21_i2_4_lut (.A(\new_sboxw[21] ), .B(n7_adj_8028), 
         .C(n33846), .D(n8_adj_8029), .Z(n2_adj_8030)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_21_i2_4_lut.init = 16'h3aca;
    LUT4 mux_692_Mux_25_i2_4_lut (.A(\round_key_gen.trw[1] ), .B(n9), .C(n33846), 
         .D(n10), .Z(n2_adj_8031)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_25_i2_4_lut.init = 16'h3aca;
    LUT4 round_key_101__bdd_3_lut_28349 (.A(round_key[101]), .B(n33846), 
         .C(\block_reg[0][5] ), .Z(n32300)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_101__bdd_3_lut_28349.init = 16'h4848;
    LUT4 \round_key_gen.trw_13__bdd_3_lut_28354  (.A(\round_key_gen.trw[13] ), 
         .B(n32302), .C(n33846), .Z(n32303)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \round_key_gen.trw_13__bdd_3_lut_28354 .init = 16'hcaca;
    LUT4 round_key_100__bdd_3_lut (.A(round_key[100]), .B(n33846), .C(\block_reg[0][4] ), 
         .Z(n32306)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_100__bdd_3_lut.init = 16'h4848;
    LUT4 \round_key_gen.trw_12__bdd_4_lut_28333  (.A(round_key[100]), .B(n28933), 
         .C(n33897), .D(n33893), .Z(n32308)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam \round_key_gen.trw_12__bdd_4_lut_28333 .init = 16'h6996;
    LUT4 \round_key_gen.trw_12__bdd_3_lut_28334  (.A(\round_key_gen.trw[12] ), 
         .B(n32308), .C(n33846), .Z(n32309)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \round_key_gen.trw_12__bdd_3_lut_28334 .init = 16'hcaca;
    LUT4 mux_692_Mux_89_i2_4_lut (.A(\round_key_gen.trw[1] ), .B(n7_adj_8032), 
         .C(n33846), .D(n8_adj_8033), .Z(n2_adj_8034)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_89_i2_4_lut.init = 16'h3aca;
    LUT4 n33038_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n33036), .D(n33038), 
         .Z(n33039)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n33038_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 round_key_96__bdd_3_lut (.A(round_key[96]), .B(n33846), .C(\block_reg[0][0] ), 
         .Z(n32321)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_96__bdd_3_lut.init = 16'h4848;
    LUT4 i4053_3_lut (.A(\enc_new_block[56] ), .B(\enc_new_block[24] ), 
         .C(n6364[3]), .Z(n9662)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam i4053_3_lut.init = 16'hcaca;
    LUT4 n33056_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n33054), .D(n33056), 
         .Z(n33057)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n33056_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n33071_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n33069), .D(n33071), 
         .Z(n33072)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n33071_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n33080_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n33078), .D(n33080), 
         .Z(n33081)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n33080_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n33092_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n33090), .D(n33092), 
         .Z(n33093)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n33092_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_178_i25_3_lut (.A(\enc_new_block[120] ), .B(\enc_new_block[88] ), 
         .C(n6364_c[1]), .Z(n2531[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam mux_178_i25_3_lut.init = 16'hcaca;
    LUT4 \round_key_gen.trw_8__bdd_4_lut_28288  (.A(round_key[96]), .B(n33897), 
         .C(n33898), .D(\enc_new_block[40] ), .Z(n32323)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam \round_key_gen.trw_8__bdd_4_lut_28288 .init = 16'h6996;
    LUT4 \round_key_gen.trw_8__bdd_3_lut_28289  (.A(\round_key_gen.trw[8] ), 
         .B(n32323), .C(n33846), .Z(n32324)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \round_key_gen.trw_8__bdd_3_lut_28289 .init = 16'hcaca;
    LUT4 round_key_95__bdd_3_lut (.A(round_key[95]), .B(n33846), .C(\block_reg[1][31] ), 
         .Z(n32327)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_95__bdd_3_lut.init = 16'h4848;
    LUT4 mux_692_Mux_91_i2_4_lut (.A(\round_key_gen.trw[3] ), .B(n7_adj_8035), 
         .C(n33846), .D(n8_adj_8036), .Z(n2_adj_8037)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_91_i2_4_lut.init = 16'h3aca;
    LUT4 i4051_3_lut (.A(\enc_new_block[55] ), .B(\enc_new_block[23] ), 
         .C(n6364[3]), .Z(n9660)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam i4051_3_lut.init = 16'hcaca;
    LUT4 n33111_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n33109), .D(n33111), 
         .Z(n33112)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n33111_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n33125_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n33123), .D(n33125), 
         .Z(n33126)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n33125_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_178_i24_3_lut (.A(\enc_new_block[119] ), .B(\enc_new_block[87] ), 
         .C(n6364_c[1]), .Z(n2531[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam mux_178_i24_3_lut.init = 16'hcaca;
    LUT4 n33134_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n33132), .D(n33134), 
         .Z(n33135)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n33134_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 \round_key_gen.trw_7__bdd_4_lut_28272  (.A(round_key[95]), .B(n33889), 
         .C(n33890), .D(\round_logic.mixcolumns_block_71__N_1149[0] ), .Z(n32329)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam \round_key_gen.trw_7__bdd_4_lut_28272 .init = 16'h6996;
    LUT4 \round_key_gen.trw_7__bdd_3_lut_28273  (.A(\round_key_gen.trw[7] ), 
         .B(n32329), .C(n33846), .Z(n32330)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \round_key_gen.trw_7__bdd_3_lut_28273 .init = 16'hcaca;
    LUT4 mux_692_Mux_92_i2_4_lut (.A(\round_key_gen.trw[4] ), .B(n7_adj_8038), 
         .C(n33846), .D(n8_adj_8039), .Z(n2_adj_8040)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_92_i2_4_lut.init = 16'h3aca;
    LUT4 i4049_3_lut (.A(\enc_new_block[54] ), .B(\enc_new_block[22] ), 
         .C(n6364[3]), .Z(n9658)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam i4049_3_lut.init = 16'hcaca;
    LUT4 round_key_94__bdd_3_lut (.A(round_key[94]), .B(n33846), .C(\block_reg[1][30] ), 
         .Z(n32333)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_94__bdd_3_lut.init = 16'h4848;
    LUT4 mux_692_Mux_27_i2_4_lut (.A(\round_key_gen.trw[3] ), .B(n7_adj_8041), 
         .C(n33846), .D(n8_adj_8042), .Z(n2_adj_8043)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_27_i2_4_lut.init = 16'h3aca;
    LUT4 mux_178_i23_3_lut (.A(\enc_new_block[118] ), .B(\enc_new_block[86] ), 
         .C(n6364_c[1]), .Z(n2531[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam mux_178_i23_3_lut.init = 16'hcaca;
    LUT4 \round_key_gen.trw_6__bdd_4_lut_28689  (.A(round_key[94]), .B(n33887), 
         .C(n33888), .D(\enc_new_block[54] ), .Z(n32335)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam \round_key_gen.trw_6__bdd_4_lut_28689 .init = 16'h6996;
    LUT4 mux_692_Mux_28_i2_4_lut (.A(\round_key_gen.trw[4] ), .B(n9_adj_8044), 
         .C(n33846), .D(n10_adj_8045), .Z(n2_adj_8046)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_28_i2_4_lut.init = 16'h3aca;
    LUT4 \round_key_gen.trw_6__bdd_3_lut_28690  (.A(\round_key_gen.trw[6] ), 
         .B(n32335), .C(n33846), .Z(n32336)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \round_key_gen.trw_6__bdd_3_lut_28690 .init = 16'hcaca;
    LUT4 mux_692_Mux_30_i2_4_lut (.A(\round_key_gen.trw[6] ), .B(n7_adj_8047), 
         .C(n33846), .D(n8_adj_8048), .Z(n2_adj_8049)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_30_i2_4_lut.init = 16'h3aca;
    LUT4 i4047_3_lut (.A(\enc_new_block[53] ), .B(\enc_new_block[21] ), 
         .C(n6364[3]), .Z(n9656)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam i4047_3_lut.init = 16'hcaca;
    LUT4 mux_178_i22_3_lut (.A(\enc_new_block[117] ), .B(\enc_new_block[85] ), 
         .C(n6364_c[1]), .Z(n2531[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam mux_178_i22_3_lut.init = 16'hcaca;
    LUT4 mux_692_Mux_33_i2_4_lut (.A(\round_key_gen.trw[9] ), .B(n7_adj_8050), 
         .C(n33846), .D(n8_adj_8051), .Z(n2_adj_8052)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_33_i2_4_lut.init = 16'h3aca;
    LUT4 mux_692_Mux_34_i2_4_lut (.A(\round_key_gen.trw[10] ), .B(n7_adj_8053), 
         .C(n33846), .D(n8_adj_8054), .Z(n2_adj_8055)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_34_i2_4_lut.init = 16'h3aca;
    LUT4 i4045_3_lut (.A(\enc_new_block[52] ), .B(\enc_new_block[20] ), 
         .C(n6364[3]), .Z(n9654)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam i4045_3_lut.init = 16'hcaca;
    LUT4 round_key_93__bdd_3_lut (.A(round_key[93]), .B(n33846), .C(\block_reg[1][29] ), 
         .Z(n32339)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_93__bdd_3_lut.init = 16'h4848;
    LUT4 mux_178_i21_3_lut (.A(\enc_new_block[116] ), .B(\enc_new_block[84] ), 
         .C(n6364_c[1]), .Z(n2531[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam mux_178_i21_3_lut.init = 16'hcaca;
    LUT4 mux_692_Mux_97_i2_4_lut (.A(\round_key_gen.trw[9] ), .B(n7_adj_8056), 
         .C(n33846), .D(n8_adj_8057), .Z(n2_adj_8058)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_97_i2_4_lut.init = 16'h3aca;
    LUT4 i4043_3_lut (.A(\enc_new_block[51] ), .B(\enc_new_block[19] ), 
         .C(n6364[3]), .Z(n9652)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam i4043_3_lut.init = 16'hcaca;
    LUT4 n33140_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n33138), .D(n33140), 
         .Z(n33141)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n33140_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 \round_key_gen.trw_5__bdd_4_lut_28823  (.A(round_key[93]), .B(n33885), 
         .C(n33886), .D(\enc_new_block[53] ), .Z(n32341)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam \round_key_gen.trw_5__bdd_4_lut_28823 .init = 16'h6996;
    LUT4 n33161_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n33159), .D(n33161), 
         .Z(n33162)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n33161_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n33175_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n33173), .D(n33175), 
         .Z(n33176)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n33175_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 \round_key_gen.trw_5__bdd_3_lut_28824  (.A(\round_key_gen.trw[5] ), 
         .B(n32341), .C(n33846), .Z(n32342)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \round_key_gen.trw_5__bdd_3_lut_28824 .init = 16'hcaca;
    LUT4 mux_178_i20_3_lut (.A(\enc_new_block[115] ), .B(\enc_new_block[83] ), 
         .C(n6364_c[1]), .Z(n2531[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam mux_178_i20_3_lut.init = 16'hcaca;
    LUT4 mux_692_Mux_98_i2_4_lut (.A(\round_key_gen.trw[10] ), .B(n7_adj_8059), 
         .C(n33846), .D(n8_adj_8060), .Z(n2_adj_8061)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_98_i2_4_lut.init = 16'h3aca;
    LUT4 mux_692_Mux_36_i2_4_lut (.A(\round_key_gen.trw[12] ), .B(n7_adj_8062), 
         .C(n33846), .D(n8_adj_8063), .Z(n2_adj_8064)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_36_i2_4_lut.init = 16'h3aca;
    LUT4 mux_692_Mux_99_i2_4_lut (.A(\round_key_gen.trw[11] ), .B(n7_adj_8065), 
         .C(n33846), .D(n8_adj_8066), .Z(n2_adj_8067)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_99_i2_4_lut.init = 16'h3aca;
    LUT4 i4041_3_lut (.A(\enc_new_block[50] ), .B(\enc_new_block[18] ), 
         .C(n6364[3]), .Z(n9650)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam i4041_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_563 (.A(\enc_new_block[58] ), .B(\enc_new_block[18] ), 
         .Z(n33867)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_rep_563.init = 16'h6666;
    LUT4 mux_692_Mux_102_i2_4_lut (.A(\round_key_gen.trw[14] ), .B(n7_adj_8068), 
         .C(n33846), .D(n8_adj_8069), .Z(n2_adj_8070)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_102_i2_4_lut.init = 16'h3aca;
    LUT4 mux_692_Mux_105_i2_4_lut (.A(\round_key_gen.trw[17] ), .B(n7_adj_8071), 
         .C(n33846), .D(n8_adj_8072), .Z(n2_adj_8073)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_105_i2_4_lut.init = 16'h3aca;
    LUT4 round_key_90__bdd_3_lut (.A(round_key[90]), .B(n33846), .C(\block_reg[1][26] ), 
         .Z(n32363)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_90__bdd_3_lut.init = 16'h4848;
    LUT4 mux_178_i19_3_lut (.A(\enc_new_block[114] ), .B(\enc_new_block[82] ), 
         .C(n6364_c[1]), .Z(n2531[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam mux_178_i19_3_lut.init = 16'hcaca;
    LUT4 n33184_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n33182), .D(n33184), 
         .Z(n33185)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n33184_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n33196_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n33194), .D(n33196), 
         .Z(n33197)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n33196_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n33208_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n33206), .D(n33208), 
         .Z(n33209)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n33208_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_692_Mux_107_i2_4_lut (.A(\round_key_gen.trw[19] ), .B(n7_adj_8074), 
         .C(n33846), .D(n8_adj_8075), .Z(n2_adj_8076)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_107_i2_4_lut.init = 16'h3aca;
    LUT4 i4039_3_lut (.A(\enc_new_block[49] ), .B(\enc_new_block[17] ), 
         .C(n6364[3]), .Z(n9648)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam i4039_3_lut.init = 16'hcaca;
    LUT4 i2_2_lut_3_lut (.A(\enc_new_block[58] ), .B(\enc_new_block[18] ), 
         .C(\enc_new_block[67] ), .Z(n7_adj_8077)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i2_2_lut_3_lut.init = 16'h9696;
    LUT4 mux_178_i18_3_lut (.A(\enc_new_block[113] ), .B(\enc_new_block[81] ), 
         .C(n6364_c[1]), .Z(n2531[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam mux_178_i18_3_lut.init = 16'hcaca;
    LUT4 mux_692_Mux_108_i2_4_lut (.A(\round_key_gen.trw[20] ), .B(n9_adj_8078), 
         .C(n33846), .D(n10_adj_8079), .Z(n2_adj_8080)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_108_i2_4_lut.init = 16'h3aca;
    LUT4 n33220_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n33218), .D(n33220), 
         .Z(n33221)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n33220_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i4037_3_lut (.A(\enc_new_block[48] ), .B(\enc_new_block[16] ), 
         .C(n6364[3]), .Z(n9646)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam i4037_3_lut.init = 16'hcaca;
    LUT4 mux_178_i17_3_lut (.A(\enc_new_block[112] ), .B(\enc_new_block[80] ), 
         .C(n6364_c[1]), .Z(n2531[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam mux_178_i17_3_lut.init = 16'hcaca;
    LUT4 i4035_3_lut (.A(\round_logic.mixcolumns_block_111__N_1285[0] ), .B(\round_logic.mixcolumns_block_79__N_1341[0] ), 
         .C(n6364[3]), .Z(n9644)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam i4035_3_lut.init = 16'hcaca;
    LUT4 mux_178_i16_3_lut (.A(\round_logic.mixcolumns_block_47__N_1397[0] ), 
         .B(\round_logic.mixcolumns_block_15__N_1453[0] ), .C(n6364_c[1]), 
         .Z(n2531[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam mux_178_i16_3_lut.init = 16'hcaca;
    LUT4 i4033_3_lut (.A(\round_logic.mixcolumns_block_111__N_1285[7] ), .B(\round_logic.mixcolumns_block_79__N_1341[7] ), 
         .C(n6364[3]), .Z(n9642)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam i4033_3_lut.init = 16'hcaca;
    LUT4 mux_178_i15_3_lut (.A(\round_logic.mixcolumns_block_47__N_1397[7] ), 
         .B(\round_logic.mixcolumns_block_15__N_1453[7] ), .C(n6364_c[1]), 
         .Z(n2531[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam mux_178_i15_3_lut.init = 16'hcaca;
    LUT4 n33226_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n33224), .D(n33226), 
         .Z(n33227)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n33226_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n33238_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n33236), .D(n33238), 
         .Z(n33239)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n33238_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_692_Mux_37_i2_4_lut (.A(\round_key_gen.trw[13] ), .B(n7_adj_8081), 
         .C(n33846), .D(n8_adj_8082), .Z(n2_adj_8083)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_37_i2_4_lut.init = 16'h3aca;
    LUT4 n33273_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n33271), .D(n33273), 
         .Z(n33274)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n33273_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_692_Mux_113_i2_4_lut (.A(\new_sboxw[17] ), .B(n7_adj_8084), 
         .C(n33846), .D(n8_adj_8085), .Z(n2_adj_8086)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_113_i2_4_lut.init = 16'h3aca;
    LUT4 i4031_3_lut (.A(\round_logic.mixcolumns_block_111__N_1285[6] ), .B(\round_logic.mixcolumns_block_79__N_1341[6] ), 
         .C(n6364[3]), .Z(n9640)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam i4031_3_lut.init = 16'hcaca;
    LUT4 mux_692_Mux_114_i2_4_lut (.A(\new_sboxw[18] ), .B(n7_adj_8087), 
         .C(n33846), .D(n8_adj_8088), .Z(n2_adj_8089)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_114_i2_4_lut.init = 16'h3aca;
    LUT4 mux_692_Mux_115_i2_4_lut (.A(\new_sboxw[19] ), .B(n7_adj_8090), 
         .C(n33846), .D(n8_adj_8091), .Z(n2_adj_8092)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_115_i2_4_lut.init = 16'h3aca;
    LUT4 mux_692_Mux_116_i2_4_lut (.A(\new_sboxw[20] ), .B(n9_adj_8093), 
         .C(n33846), .D(n10_adj_8094), .Z(n2_adj_8095)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_116_i2_4_lut.init = 16'h3aca;
    LUT4 mux_692_Mux_39_i2_4_lut (.A(\round_key_gen.trw[15] ), .B(n7_adj_8096), 
         .C(n33846), .D(n8_adj_8097), .Z(n2_adj_8098)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_39_i2_4_lut.init = 16'h3aca;
    LUT4 mux_692_Mux_118_i2_4_lut (.A(\new_sboxw[22] ), .B(n7_adj_8099), 
         .C(n33846), .D(n8_adj_8100), .Z(n2_adj_8101)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_118_i2_4_lut.init = 16'h3aca;
    LUT4 mux_692_Mux_119_i2_4_lut (.A(\new_sboxw[23] ), .B(n7_adj_8102), 
         .C(n33846), .D(n8_adj_8103), .Z(n2_adj_8104)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_119_i2_4_lut.init = 16'h3aca;
    LUT4 i3_3_lut_4_lut (.A(\enc_new_block[58] ), .B(\enc_new_block[18] ), 
         .C(\enc_new_block[57] ), .D(\round_logic.mixcolumns_block_39__N_1197[2] ), 
         .Z(n8_adj_8054)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i3_3_lut_4_lut.init = 16'h6996;
    LUT4 mux_692_Mux_41_i2_4_lut (.A(\round_key_gen.trw[17] ), .B(n7_adj_8105), 
         .C(n33846), .D(n8_adj_8106), .Z(n2_adj_8107)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_41_i2_4_lut.init = 16'h3aca;
    LUT4 mux_692_Mux_121_i2_4_lut (.A(\round_key_gen.trw[1] ), .B(n7_adj_8108), 
         .C(n33846), .D(n8_adj_8109), .Z(n2_adj_8110)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_121_i2_4_lut.init = 16'h3aca;
    LUT4 mux_692_Mux_123_i2_4_lut (.A(\round_key_gen.trw[3] ), .B(n7_adj_8111), 
         .C(n33846), .D(n8_adj_8112), .Z(n2_adj_8113)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_123_i2_4_lut.init = 16'h3aca;
    LUT4 mux_692_Mux_125_i2_4_lut (.A(\round_key_gen.trw[5] ), .B(n7_adj_8114), 
         .C(n33846), .D(n8_adj_8115), .Z(n2_adj_8116)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_125_i2_4_lut.init = 16'h3aca;
    PFUMX i28975 (.BLUT(n33270), .ALUT(n33269), .C0(n33847), .Z(n33271));
    LUT4 mux_178_i14_3_lut (.A(\round_logic.mixcolumns_block_47__N_1397[6] ), 
         .B(\round_logic.mixcolumns_block_15__N_1453[6] ), .C(n6364_c[1]), 
         .Z(n2531[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam mux_178_i14_3_lut.init = 16'hcaca;
    LUT4 mux_692_Mux_43_i2_4_lut (.A(\round_key_gen.trw[19] ), .B(n7_adj_8117), 
         .C(n33846), .D(n8_adj_8118), .Z(n2_adj_8119)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_43_i2_4_lut.init = 16'h3aca;
    LUT4 i4029_3_lut (.A(\round_logic.mixcolumns_block_111__N_1285[5] ), .B(\round_logic.mixcolumns_block_79__N_1341[5] ), 
         .C(n6364[3]), .Z(n9638)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam i4029_3_lut.init = 16'hcaca;
    LUT4 round_key_0__bdd_3_lut_28974_4_lut_4_lut (.A(n33846), .B(round_key[0]), 
         .C(\enc_new_block[32] ), .D(n33845), .Z(n33269)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_0__bdd_3_lut_28974_4_lut_4_lut.init = 16'h1400;
    LUT4 round_key_6__bdd_3_lut_28944_4_lut_4_lut (.A(n33846), .B(round_key[6]), 
         .C(\round_logic.mixcolumns_block_7__N_1245[7] ), .D(n33845), .Z(n33234)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_6__bdd_3_lut_28944_4_lut_4_lut.init = 16'h1400;
    LUT4 mux_178_i13_3_lut (.A(\round_logic.mixcolumns_block_47__N_1397[5] ), 
         .B(\round_logic.mixcolumns_block_15__N_1453[5] ), .C(n6364_c[1]), 
         .Z(n2531[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam mux_178_i13_3_lut.init = 16'hcaca;
    LUT4 i4027_3_lut (.A(\enc_new_block[43] ), .B(\enc_new_block[11] ), 
         .C(n6364[3]), .Z(n9636)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam i4027_3_lut.init = 16'hcaca;
    LUT4 mux_178_i12_3_lut (.A(\enc_new_block[107] ), .B(\enc_new_block[75] ), 
         .C(n6364_c[1]), .Z(n2531[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam mux_178_i12_3_lut.init = 16'hcaca;
    LUT4 round_key_8__bdd_3_lut_28933_4_lut_4_lut (.A(n33846), .B(round_key[8]), 
         .C(\enc_new_block[72] ), .D(n33845), .Z(n33222)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_8__bdd_3_lut_28933_4_lut_4_lut.init = 16'h1400;
    LUT4 \round_key_gen.trw_2__bdd_4_lut_28648  (.A(round_key[90]), .B(n33878), 
         .C(n33879), .D(\enc_new_block[50] ), .Z(n32365)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam \round_key_gen.trw_2__bdd_4_lut_28648 .init = 16'h6996;
    LUT4 round_key_9__bdd_3_lut_28930_4_lut_4_lut (.A(n33846), .B(round_key[9]), 
         .C(\round_logic.mixcolumns_block_15__N_1453[2] ), .D(n33845), .Z(n33216)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_9__bdd_3_lut_28930_4_lut_4_lut.init = 16'h1400;
    LUT4 round_key_11__bdd_3_lut_28920_4_lut_4_lut (.A(n33846), .B(round_key[11]), 
         .C(\enc_new_block[75] ), .D(n33845), .Z(n33204)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_11__bdd_3_lut_28920_4_lut_4_lut.init = 16'h1400;
    LUT4 round_key_13__bdd_3_lut_28910_4_lut_4_lut (.A(n33846), .B(round_key[13]), 
         .C(\round_logic.mixcolumns_block_15__N_1453[6] ), .D(n33845), .Z(n33192)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_13__bdd_3_lut_28910_4_lut_4_lut.init = 16'h1400;
    LUT4 i4025_3_lut (.A(\enc_new_block[42] ), .B(\enc_new_block[10] ), 
         .C(n6364[3]), .Z(n9634)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam i4025_3_lut.init = 16'hcaca;
    LUT4 round_key_15__bdd_3_lut_28899_4_lut_4_lut (.A(n33846), .B(round_key[15]), 
         .C(\round_logic.mixcolumns_block_15__N_1453[0] ), .D(n33845), .Z(n33180)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_15__bdd_3_lut_28899_4_lut_4_lut.init = 16'h1400;
    LUT4 round_key_16__bdd_3_lut_28891_4_lut_4_lut (.A(n33846), .B(round_key[16]), 
         .C(\enc_new_block[112] ), .D(n33845), .Z(n33171)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_16__bdd_3_lut_28891_4_lut_4_lut.init = 16'h1400;
    LUT4 mux_178_i11_3_lut (.A(\enc_new_block[106] ), .B(\enc_new_block[74] ), 
         .C(n6364_c[1]), .Z(n2531[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam mux_178_i11_3_lut.init = 16'hcaca;
    LUT4 round_key_18__bdd_3_lut_28881_4_lut_4_lut (.A(n33846), .B(round_key[18]), 
         .C(\enc_new_block[114] ), .D(n33845), .Z(n33157)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_18__bdd_3_lut_28881_4_lut_4_lut.init = 16'h1400;
    LUT4 round_key_22__bdd_3_lut_28861_4_lut_4_lut (.A(n33846), .B(round_key[22]), 
         .C(\enc_new_block[118] ), .D(n33845), .Z(n33136)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_22__bdd_3_lut_28861_4_lut_4_lut.init = 16'h1400;
    LUT4 i4023_3_lut (.A(\round_logic.mixcolumns_block_111__N_1285[2] ), .B(\round_logic.mixcolumns_block_79__N_1341[2] ), 
         .C(n6364[3]), .Z(n9632)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam i4023_3_lut.init = 16'hcaca;
    LUT4 mux_692_Mux_44_i2_4_lut (.A(\round_key_gen.trw[20] ), .B(n7_adj_8120), 
         .C(n33846), .D(n8_adj_8121), .Z(n2_adj_8122)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_44_i2_4_lut.init = 16'h3aca;
    LUT4 mux_178_i10_3_lut (.A(\round_logic.mixcolumns_block_47__N_1397[2] ), 
         .B(\round_logic.mixcolumns_block_15__N_1453[2] ), .C(n6364_c[1]), 
         .Z(n2531[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam mux_178_i10_3_lut.init = 16'hcaca;
    LUT4 round_key_23__bdd_3_lut_28856_4_lut_4_lut (.A(n33846), .B(round_key[23]), 
         .C(\enc_new_block[119] ), .D(n33845), .Z(n33130)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_23__bdd_3_lut_28856_4_lut_4_lut.init = 16'h1400;
    LUT4 \round_key_gen.trw_2__bdd_3_lut_28649  (.A(\round_key_gen.trw[2] ), 
         .B(n32365), .C(n33846), .Z(n32366)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \round_key_gen.trw_2__bdd_3_lut_28649 .init = 16'hcaca;
    LUT4 round_key_24__bdd_3_lut_28848_4_lut_4_lut (.A(n33846), .B(round_key[24]), 
         .C(\enc_new_block[24] ), .D(n33845), .Z(n33121)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_24__bdd_3_lut_28848_4_lut_4_lut.init = 16'h1400;
    LUT4 round_key_26__bdd_3_lut_28836_4_lut_4_lut (.A(n33846), .B(round_key[26]), 
         .C(\enc_new_block[26] ), .D(n33845), .Z(n33107)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_26__bdd_3_lut_28836_4_lut_4_lut.init = 16'h1400;
    LUT4 i4021_3_lut (.A(\enc_new_block[40] ), .B(\enc_new_block[8] ), .C(n6364[3]), 
         .Z(n9630)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam i4021_3_lut.init = 16'hcaca;
    LUT4 mux_178_i9_3_lut (.A(\enc_new_block[104] ), .B(\enc_new_block[72] ), 
         .C(n6364_c[1]), .Z(n2531[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam mux_178_i9_3_lut.init = 16'hcaca;
    LUT4 round_key_29__bdd_3_lut_28820_4_lut_4_lut (.A(n33846), .B(round_key[29]), 
         .C(\enc_new_block[29] ), .D(n33845), .Z(n33088)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_29__bdd_3_lut_28820_4_lut_4_lut.init = 16'h1400;
    LUT4 i4019_3_lut (.A(\round_logic.mixcolumns_block_7__N_1245[0] ), .B(\round_logic.mixcolumns_block_103__N_1101[0] ), 
         .C(n6364[3]), .Z(n9628)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam i4019_3_lut.init = 16'hcaca;
    LUT4 round_key_31__bdd_3_lut_28811_4_lut_4_lut (.A(n33846), .B(round_key[31]), 
         .C(\enc_new_block[31] ), .D(n33845), .Z(n33076)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_31__bdd_3_lut_28811_4_lut_4_lut.init = 16'h1400;
    LUT4 round_key_32__bdd_3_lut_28805_4_lut_4_lut (.A(n33846), .B(round_key[32]), 
         .C(\enc_new_block[64] ), .D(n33845), .Z(n33067)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_32__bdd_3_lut_28805_4_lut_4_lut.init = 16'h1400;
    LUT4 round_key_35__bdd_3_lut_28792_4_lut_4_lut (.A(n33846), .B(round_key[35]), 
         .C(\enc_new_block[67] ), .D(n33845), .Z(n33052)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_35__bdd_3_lut_28792_4_lut_4_lut.init = 16'h1400;
    LUT4 mux_178_i8_3_lut (.A(\round_logic.mixcolumns_block_71__N_1149[0] ), 
         .B(\round_logic.mixcolumns_block_39__N_1197[0] ), .C(n6364_c[1]), 
         .Z(n2531[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam mux_178_i8_3_lut.init = 16'hcaca;
    LUT4 round_key_38__bdd_3_lut_28777_4_lut_4_lut (.A(n33846), .B(round_key[38]), 
         .C(\round_logic.mixcolumns_block_39__N_1197[7] ), .D(n33845), .Z(n33034)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_38__bdd_3_lut_28777_4_lut_4_lut.init = 16'h1400;
    LUT4 i4017_3_lut (.A(\round_logic.mixcolumns_block_7__N_1245[7] ), .B(\round_logic.mixcolumns_block_103__N_1101[7] ), 
         .C(n6364[3]), .Z(n9626)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam i4017_3_lut.init = 16'hcaca;
    LUT4 mux_178_i7_3_lut (.A(\round_logic.mixcolumns_block_71__N_1149[7] ), 
         .B(\round_logic.mixcolumns_block_39__N_1197[7] ), .C(n6364_c[1]), 
         .Z(n2531[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam mux_178_i7_3_lut.init = 16'hcaca;
    LUT4 \round_key_gen.trw_11__bdd_3_lut_28795_4_lut  (.A(\enc_new_block[107] ), 
         .B(\enc_new_block[19] ), .C(n10_adj_8123), .D(round_key[35]), 
         .Z(n33055)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam \round_key_gen.trw_11__bdd_3_lut_28795_4_lut .init = 16'h6996;
    LUT4 round_key_40__bdd_3_lut_28766_4_lut_4_lut (.A(n33846), .B(round_key[40]), 
         .C(\enc_new_block[104] ), .D(n33845), .Z(n33022)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_40__bdd_3_lut_28766_4_lut_4_lut.init = 16'h1400;
    LUT4 i4015_3_lut (.A(\round_logic.mixcolumns_block_7__N_1245[6] ), .B(\round_logic.mixcolumns_block_103__N_1101[6] ), 
         .C(n6364[3]), .Z(n9624)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam i4015_3_lut.init = 16'hcaca;
    LUT4 mux_178_i6_3_lut (.A(\round_logic.mixcolumns_block_71__N_1149[6] ), 
         .B(\round_logic.mixcolumns_block_39__N_1197[6] ), .C(n6364_c[1]), 
         .Z(n2531[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam mux_178_i6_3_lut.init = 16'hcaca;
    LUT4 round_key_42__bdd_3_lut_28757_4_lut_4_lut (.A(n33846), .B(round_key[42]), 
         .C(\enc_new_block[106] ), .D(n33845), .Z(n33010)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_42__bdd_3_lut_28757_4_lut_4_lut.init = 16'h1400;
    LUT4 round_key_45__bdd_3_lut_28743_4_lut_4_lut (.A(n33846), .B(round_key[45]), 
         .C(\round_logic.mixcolumns_block_47__N_1397[6] ), .D(n33845), .Z(n32993)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_45__bdd_3_lut_28743_4_lut_4_lut.init = 16'h1400;
    LUT4 i4013_3_lut (.A(\round_logic.mixcolumns_block_7__N_1245[5] ), .B(\round_logic.mixcolumns_block_103__N_1101[5] ), 
         .C(n6364[3]), .Z(n9622)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam i4013_3_lut.init = 16'hcaca;
    LUT4 mux_178_i5_3_lut (.A(\round_logic.mixcolumns_block_71__N_1149[5] ), 
         .B(\round_logic.mixcolumns_block_39__N_1197[5] ), .C(n6364_c[1]), 
         .Z(n2531[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam mux_178_i5_3_lut.init = 16'hcaca;
    LUT4 round_key_46__bdd_3_lut_28737_4_lut_4_lut (.A(n33846), .B(round_key[46]), 
         .C(\round_logic.mixcolumns_block_47__N_1397[7] ), .D(n33845), .Z(n32984)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_46__bdd_3_lut_28737_4_lut_4_lut.init = 16'h1400;
    LUT4 i4011_3_lut (.A(\enc_new_block[35] ), .B(\enc_new_block[3] ), .C(n6364[3]), 
         .Z(n9620)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam i4011_3_lut.init = 16'hcaca;
    LUT4 mux_178_i4_3_lut (.A(\enc_new_block[99] ), .B(\enc_new_block[67] ), 
         .C(n6364_c[1]), .Z(n2531[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam mux_178_i4_3_lut.init = 16'hcaca;
    LUT4 round_key_47__bdd_3_lut_28734_4_lut_4_lut (.A(n33846), .B(round_key[47]), 
         .C(\round_logic.mixcolumns_block_47__N_1397[0] ), .D(n33845), .Z(n32978)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_47__bdd_3_lut_28734_4_lut_4_lut.init = 16'h1400;
    LUT4 i4009_3_lut (.A(\enc_new_block[34] ), .B(\enc_new_block[2] ), .C(n6364[3]), 
         .Z(n9618)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam i4009_3_lut.init = 16'hcaca;
    LUT4 round_key_48__bdd_3_lut_28728_4_lut_4_lut (.A(n33846), .B(round_key[48]), 
         .C(\enc_new_block[16] ), .D(n33845), .Z(n32969)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_48__bdd_3_lut_28728_4_lut_4_lut.init = 16'h1400;
    LUT4 mux_178_i3_3_lut (.A(\enc_new_block[98] ), .B(\enc_new_block[66] ), 
         .C(n6364_c[1]), .Z(n2531[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam mux_178_i3_3_lut.init = 16'hcaca;
    LUT4 round_key_52__bdd_3_lut_28710_4_lut_4_lut (.A(n33846), .B(round_key[52]), 
         .C(\enc_new_block[20] ), .D(n33845), .Z(n32948)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_52__bdd_3_lut_28710_4_lut_4_lut.init = 16'h1400;
    LUT4 round_key_53__bdd_3_lut_28704_4_lut_4_lut (.A(n33846), .B(round_key[53]), 
         .C(\enc_new_block[21] ), .D(n33845), .Z(n32939)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_53__bdd_3_lut_28704_4_lut_4_lut.init = 16'h1400;
    LUT4 round_key_54__bdd_3_lut_28701_4_lut_4_lut (.A(n33846), .B(round_key[54]), 
         .C(\enc_new_block[22] ), .D(n33845), .Z(n32933)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_54__bdd_3_lut_28701_4_lut_4_lut.init = 16'h1400;
    LUT4 i3_3_lut_4_lut_adj_331 (.A(\enc_new_block[107] ), .B(\enc_new_block[19] ), 
         .C(round_key[59]), .D(n33868), .Z(n8_adj_8124)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i3_3_lut_4_lut_adj_331.init = 16'h6996;
    LUT4 round_key_55__bdd_3_lut_28691_4_lut_4_lut (.A(n33846), .B(round_key[55]), 
         .C(\enc_new_block[23] ), .D(n33845), .Z(n32919)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_55__bdd_3_lut_28691_4_lut_4_lut.init = 16'h1400;
    LUT4 i4007_3_lut (.A(\round_logic.mixcolumns_block_7__N_1245[2] ), .B(\round_logic.mixcolumns_block_103__N_1101[2] ), 
         .C(n6364[3]), .Z(n9616)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam i4007_3_lut.init = 16'hcaca;
    LUT4 round_key_56__bdd_3_lut_28684_4_lut_4_lut (.A(n33846), .B(round_key[56]), 
         .C(\enc_new_block[56] ), .D(n33845), .Z(n32909)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_56__bdd_3_lut_28684_4_lut_4_lut.init = 16'h1400;
    LUT4 round_key_58__bdd_3_lut_28675_4_lut_4_lut (.A(n33846), .B(round_key[58]), 
         .C(\enc_new_block[58] ), .D(n33845), .Z(n32896)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_58__bdd_3_lut_28675_4_lut_4_lut.init = 16'h1400;
    LUT4 round_key_63__bdd_3_lut_28637_4_lut_4_lut (.A(n33846), .B(round_key[63]), 
         .C(\enc_new_block[63] ), .D(n33845), .Z(n32850)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_63__bdd_3_lut_28637_4_lut_4_lut.init = 16'h1400;
    LUT4 mux_178_i2_3_lut (.A(\round_logic.mixcolumns_block_71__N_1149[2] ), 
         .B(\round_logic.mixcolumns_block_39__N_1197[2] ), .C(n6364_c[1]), 
         .Z(n2531[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam mux_178_i2_3_lut.init = 16'hcaca;
    LUT4 round_key_66__bdd_3_lut_28588_4_lut_4_lut (.A(n33846), .B(round_key[66]), 
         .C(\enc_new_block[98] ), .D(n33845), .Z(n32784)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_66__bdd_3_lut_28588_4_lut_4_lut.init = 16'h1400;
    LUT4 round_key_72__bdd_3_lut_28522_4_lut_4_lut (.A(n33846), .B(round_key[72]), 
         .C(\enc_new_block[8] ), .D(n33845), .Z(n32697)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_72__bdd_3_lut_28522_4_lut_4_lut.init = 16'h1400;
    LUT4 round_key_74__bdd_3_lut_28445_4_lut_4_lut (.A(n33846), .B(round_key[74]), 
         .C(\enc_new_block[10] ), .D(n33845), .Z(n32600)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_74__bdd_3_lut_28445_4_lut_4_lut.init = 16'h1400;
    LUT4 round_key_77__bdd_3_lut_28425_4_lut_4_lut (.A(n33846), .B(round_key[77]), 
         .C(\round_logic.mixcolumns_block_79__N_1341[6] ), .D(n33845), .Z(n32577)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_77__bdd_3_lut_28425_4_lut_4_lut.init = 16'h1400;
    LUT4 i3091_3_lut (.A(\enc_new_block[32] ), .B(\enc_new_block[0] ), .C(n6364[3]), 
         .Z(n8532)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam i3091_3_lut.init = 16'hcaca;
    LUT4 round_key_78__bdd_3_lut_28420_4_lut_4_lut (.A(n33846), .B(round_key[78]), 
         .C(\round_logic.mixcolumns_block_79__N_1341[7] ), .D(n33845), .Z(n32571)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_78__bdd_3_lut_28420_4_lut_4_lut.init = 16'h1400;
    LUT4 round_key_79__bdd_3_lut_28412_4_lut_4_lut (.A(n33846), .B(round_key[79]), 
         .C(\round_logic.mixcolumns_block_79__N_1341[0] ), .D(n33845), .Z(n32560)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_79__bdd_3_lut_28412_4_lut_4_lut.init = 16'h1400;
    LUT4 round_key_80__bdd_3_lut_28407_4_lut_4_lut (.A(n33846), .B(round_key[80]), 
         .C(\enc_new_block[48] ), .D(n33845), .Z(n32554)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_80__bdd_3_lut_28407_4_lut_4_lut.init = 16'h1400;
    LUT4 mux_178_i1_3_lut (.A(\enc_new_block[96] ), .B(\enc_new_block[64] ), 
         .C(n6364_c[1]), .Z(n2531[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam mux_178_i1_3_lut.init = 16'hcaca;
    LUT4 round_key_88__bdd_3_lut_28368_4_lut_4_lut (.A(n33846), .B(round_key[88]), 
         .C(\enc_new_block[88] ), .D(n33845), .Z(n32508)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_88__bdd_3_lut_28368_4_lut_4_lut.init = 16'h1400;
    LUT4 round_key_90__bdd_3_lut_28281_4_lut_4_lut (.A(n33846), .B(round_key[90]), 
         .C(\enc_new_block[90] ), .D(n33845), .Z(n32362)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_90__bdd_3_lut_28281_4_lut_4_lut.init = 16'h1400;
    LUT4 round_key_93__bdd_3_lut_28264_4_lut_4_lut (.A(n33846), .B(round_key[93]), 
         .C(\enc_new_block[93] ), .D(n33845), .Z(n32338)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_93__bdd_3_lut_28264_4_lut_4_lut.init = 16'h1400;
    LUT4 round_key_94__bdd_3_lut_28259_4_lut_4_lut (.A(n33846), .B(round_key[94]), 
         .C(\enc_new_block[94] ), .D(n33845), .Z(n32332)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_94__bdd_3_lut_28259_4_lut_4_lut.init = 16'h1400;
    LUT4 round_key_95__bdd_3_lut_28254_4_lut_4_lut (.A(n33846), .B(round_key[95]), 
         .C(\enc_new_block[95] ), .D(n33845), .Z(n32326)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_95__bdd_3_lut_28254_4_lut_4_lut.init = 16'h1400;
    LUT4 round_key_96__bdd_3_lut_28251_4_lut_4_lut (.A(n33846), .B(round_key[96]), 
         .C(\enc_new_block[0] ), .D(n33845), .Z(n32320)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_96__bdd_3_lut_28251_4_lut_4_lut.init = 16'h1400;
    LUT4 round_key_100__bdd_3_lut_28239_4_lut_4_lut (.A(n33846), .B(round_key[100]), 
         .C(\round_logic.mixcolumns_block_103__N_1101[5] ), .D(n33845), 
         .Z(n32305)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_100__bdd_3_lut_28239_4_lut_4_lut.init = 16'h1400;
    LUT4 round_key_101__bdd_3_lut_28235_4_lut_4_lut (.A(n33846), .B(round_key[101]), 
         .C(\round_logic.mixcolumns_block_103__N_1101[6] ), .D(n33845), 
         .Z(n32299)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_101__bdd_3_lut_28235_4_lut_4_lut.init = 16'h1400;
    LUT4 round_key_103__bdd_3_lut_28229_4_lut_4_lut (.A(n33846), .B(round_key[103]), 
         .C(\round_logic.mixcolumns_block_103__N_1101[0] ), .D(n33845), 
         .Z(n32290)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_103__bdd_3_lut_28229_4_lut_4_lut.init = 16'h1400;
    LUT4 round_key_104__bdd_3_lut_28225_4_lut_4_lut (.A(n33846), .B(round_key[104]), 
         .C(\enc_new_block[40] ), .D(n33845), .Z(n32284)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_104__bdd_3_lut_28225_4_lut_4_lut.init = 16'h1400;
    LUT4 round_key_106__bdd_3_lut_28219_4_lut_4_lut (.A(n33846), .B(round_key[106]), 
         .C(\enc_new_block[42] ), .D(n33845), .Z(n32275)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_106__bdd_3_lut_28219_4_lut_4_lut.init = 16'h1400;
    LUT4 round_key_109__bdd_3_lut_28209_4_lut_4_lut (.A(n33846), .B(round_key[109]), 
         .C(\round_logic.mixcolumns_block_111__N_1285[6] ), .D(n33845), 
         .Z(n32261)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_109__bdd_3_lut_28209_4_lut_4_lut.init = 16'h1400;
    LUT4 round_key_110__bdd_3_lut_28206_4_lut_4_lut (.A(n33846), .B(round_key[110]), 
         .C(\round_logic.mixcolumns_block_111__N_1285[7] ), .D(n33845), 
         .Z(n32255)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_110__bdd_3_lut_28206_4_lut_4_lut.init = 16'h1400;
    LUT4 round_key_111__bdd_3_lut_28203_4_lut_4_lut (.A(n33846), .B(round_key[111]), 
         .C(\round_logic.mixcolumns_block_111__N_1285[0] ), .D(n33845), 
         .Z(n32249)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_111__bdd_3_lut_28203_4_lut_4_lut.init = 16'h1400;
    LUT4 round_key_112__bdd_3_lut_28200_4_lut_4_lut (.A(n33846), .B(round_key[112]), 
         .C(\enc_new_block[80] ), .D(n33845), .Z(n32243)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_112__bdd_3_lut_28200_4_lut_4_lut.init = 16'h1400;
    LUT4 round_key_117__bdd_3_lut_28184_4_lut_4_lut (.A(n33846), .B(round_key[117]), 
         .C(\enc_new_block[85] ), .D(n33845), .Z(n32223)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_117__bdd_3_lut_28184_4_lut_4_lut.init = 16'h1400;
    LUT4 round_key_120__bdd_3_lut_28175_4_lut_4_lut (.A(n33846), .B(round_key[120]), 
         .C(\enc_new_block[120] ), .D(n33845), .Z(n32211)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_120__bdd_3_lut_28175_4_lut_4_lut.init = 16'h1400;
    LUT4 round_key_122__bdd_3_lut_28169_4_lut_4_lut (.A(n33846), .B(round_key[122]), 
         .C(\enc_new_block[122] ), .D(n33845), .Z(n32202)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_122__bdd_3_lut_28169_4_lut_4_lut.init = 16'h1400;
    LUT4 i15389_3_lut_4_lut_4_lut (.A(n33846), .B(\enc_new_block[27] ), 
         .C(round_key[27]), .D(n33845), .Z(n12960)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i15389_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i15388_3_lut_4_lut_4_lut (.A(n33846), .B(\enc_new_block[28] ), 
         .C(round_key[28]), .D(n33845), .Z(n12961)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i15388_3_lut_4_lut_4_lut.init = 16'h1400;
    FD1P3AX block_w3_reg__i1 (.D(n33274), .SP(block_w3_we), .CK(clk_c), 
            .Q(\enc_new_block[0] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w3_reg__i1.GSR = "ENABLED";
    LUT4 i15386_3_lut_4_lut_4_lut (.A(n33846), .B(\enc_new_block[30] ), 
         .C(round_key[30]), .D(n33845), .Z(n12963)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i15386_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i15383_3_lut_4_lut_4_lut (.A(n33846), .B(\round_logic.mixcolumns_block_39__N_1197[2] ), 
         .C(round_key[33]), .D(n33845), .Z(n12966)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i15383_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i15382_3_lut_4_lut_4_lut (.A(n33846), .B(\enc_new_block[66] ), 
         .C(round_key[34]), .D(n33845), .Z(n12967)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i15382_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i15419_3_lut_4_lut_4_lut (.A(n33846), .B(\round_logic.mixcolumns_block_39__N_1197[5] ), 
         .C(round_key[36]), .D(n33845), .Z(n12969)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i15419_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i14569_3_lut_4_lut_4_lut (.A(n33846), .B(\round_logic.mixcolumns_block_39__N_1197[6] ), 
         .C(round_key[37]), .D(n33845), .Z(n12970)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14569_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i14567_3_lut_4_lut_4_lut (.A(n33846), .B(\round_logic.mixcolumns_block_39__N_1197[0] ), 
         .C(round_key[39]), .D(n33845), .Z(n12972)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14567_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 mux_692_Mux_49_i2_4_lut (.A(\new_sboxw[17] ), .B(n7_adj_8125), 
         .C(n33846), .D(n8_adj_8126), .Z(n2_adj_8127)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_49_i2_4_lut.init = 16'h3aca;
    LUT4 i14565_3_lut_4_lut_4_lut (.A(n33846), .B(\round_logic.mixcolumns_block_47__N_1397[2] ), 
         .C(round_key[41]), .D(n33845), .Z(n12974)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14565_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i14563_3_lut_4_lut_4_lut (.A(n33846), .B(\enc_new_block[107] ), 
         .C(round_key[43]), .D(n33845), .Z(n12976)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14563_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i14562_3_lut_4_lut_4_lut (.A(n33846), .B(\round_logic.mixcolumns_block_47__N_1397[5] ), 
         .C(round_key[44]), .D(n33845), .Z(n12977)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14562_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 mux_692_Mux_50_i2_4_lut (.A(\new_sboxw[18] ), .B(n7_adj_8128), 
         .C(n33846), .D(n8_adj_8129), .Z(n2_adj_8130)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_50_i2_4_lut.init = 16'h3aca;
    LUT4 mux_692_Mux_51_i2_4_lut (.A(\new_sboxw[19] ), .B(n7_adj_8131), 
         .C(n33846), .D(n8_adj_8132), .Z(n2_adj_8133)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_51_i2_4_lut.init = 16'h3aca;
    LUT4 i14557_3_lut_4_lut_4_lut (.A(n33846), .B(\enc_new_block[17] ), 
         .C(round_key[49]), .D(n33845), .Z(n12982)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14557_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i14556_3_lut_4_lut_4_lut (.A(n33846), .B(\enc_new_block[18] ), 
         .C(round_key[50]), .D(n33845), .Z(n12983)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14556_3_lut_4_lut_4_lut.init = 16'h1400;
    PFUMX i28945 (.BLUT(n33235), .ALUT(n33234), .C0(n33847), .Z(n33236));
    LUT4 i14555_3_lut_4_lut_4_lut (.A(n33846), .B(\enc_new_block[19] ), 
         .C(round_key[51]), .D(n33845), .Z(n12984)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14555_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i14549_3_lut_4_lut_4_lut (.A(n33846), .B(\enc_new_block[57] ), 
         .C(round_key[57]), .D(n33845), .Z(n12990)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14549_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i1_2_lut_rep_564 (.A(\enc_new_block[23] ), .B(\enc_new_block[63] ), 
         .Z(n33868)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_rep_564.init = 16'h6666;
    LUT4 round_key_127__bdd_3_lut (.A(round_key[127]), .B(n33846), .C(\block_reg[0][31] ), 
         .Z(n32177)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_127__bdd_3_lut.init = 16'h4848;
    LUT4 \round_key_gen.trw_7__bdd_4_lut_28257  (.A(round_key[127]), .B(n29399), 
         .C(n33908), .D(\round_logic.mixcolumns_block_111__N_1285[0] ), 
         .Z(n32179)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam \round_key_gen.trw_7__bdd_4_lut_28257 .init = 16'h6996;
    LUT4 \round_key_gen.trw_7__bdd_3_lut_28258  (.A(\round_key_gen.trw[7] ), 
         .B(n32179), .C(n33846), .Z(n32180)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \round_key_gen.trw_7__bdd_3_lut_28258 .init = 16'hcaca;
    FD1P3AX block_w0_reg__i1 (.D(n32325), .SP(block_w0_we), .CK(clk_c), 
            .Q(\enc_new_block[96] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w0_reg__i1.GSR = "ENABLED";
    LUT4 i14547_3_lut_4_lut_4_lut (.A(n33846), .B(\enc_new_block[59] ), 
         .C(round_key[59]), .D(n33845), .Z(n12992)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14547_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i14546_3_lut_4_lut_4_lut (.A(n33846), .B(\enc_new_block[60] ), 
         .C(round_key[60]), .D(n33845), .Z(n12993)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14546_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i14545_3_lut_4_lut_4_lut (.A(n33846), .B(\enc_new_block[61] ), 
         .C(round_key[61]), .D(n33845), .Z(n12994)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14545_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i14544_3_lut_4_lut_4_lut (.A(n33846), .B(\enc_new_block[62] ), 
         .C(round_key[62]), .D(n33845), .Z(n12995)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14544_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 round_key_126__bdd_3_lut (.A(round_key[126]), .B(n33846), .C(\block_reg[0][30] ), 
         .Z(n32183)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_126__bdd_3_lut.init = 16'h4848;
    LUT4 i14542_3_lut_4_lut_4_lut (.A(n33846), .B(\enc_new_block[96] ), 
         .C(round_key[64]), .D(n33845), .Z(n12997)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14542_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i14541_3_lut_4_lut_4_lut (.A(n33846), .B(\round_logic.mixcolumns_block_71__N_1149[2] ), 
         .C(round_key[65]), .D(n33845), .Z(n12998)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14541_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i14539_3_lut_4_lut_4_lut (.A(n33846), .B(\enc_new_block[99] ), 
         .C(round_key[67]), .D(n33845), .Z(n13000)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14539_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i14538_3_lut_4_lut_4_lut (.A(n33846), .B(\round_logic.mixcolumns_block_71__N_1149[5] ), 
         .C(round_key[68]), .D(n33845), .Z(n13001)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14538_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 \round_key_gen.trw_6__bdd_4_lut_28262  (.A(round_key[126]), .B(n33906), 
         .C(n33907), .D(\enc_new_block[86] ), .Z(n32185)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam \round_key_gen.trw_6__bdd_4_lut_28262 .init = 16'h6996;
    LUT4 i14537_3_lut_4_lut_4_lut (.A(n33846), .B(\round_logic.mixcolumns_block_71__N_1149[6] ), 
         .C(round_key[69]), .D(n33845), .Z(n13002)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14537_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 \round_key_gen.trw_6__bdd_3_lut_28263  (.A(\round_key_gen.trw[6] ), 
         .B(n32185), .C(n33846), .Z(n32186)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \round_key_gen.trw_6__bdd_3_lut_28263 .init = 16'hcaca;
    LUT4 mux_692_Mux_57_i2_4_lut (.A(\round_key_gen.trw[1] ), .B(n7_adj_8134), 
         .C(n33846), .D(n8_adj_8135), .Z(n2_adj_8136)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_57_i2_4_lut.init = 16'h3aca;
    PFUMX i28934 (.BLUT(n33223), .ALUT(n33222), .C0(n33847), .Z(n33224));
    LUT4 i3_3_lut_4_lut_adj_332 (.A(\enc_new_block[23] ), .B(\enc_new_block[63] ), 
         .C(\enc_new_block[59] ), .D(n28939), .Z(n8_adj_8137)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i3_3_lut_4_lut_adj_332.init = 16'h6996;
    LUT4 round_key_124__bdd_3_lut (.A(round_key[124]), .B(n33846), .C(\block_reg[0][28] ), 
         .Z(n32194)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_124__bdd_3_lut.init = 16'h4848;
    LUT4 mux_692_Mux_59_i2_4_lut (.A(\round_key_gen.trw[3] ), .B(n7_adj_8077), 
         .C(n33846), .D(n8_adj_8124), .Z(n2_adj_8138)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_59_i2_4_lut.init = 16'h3aca;
    LUT4 \round_key_gen.trw_4__bdd_4_lut_28661  (.A(round_key[124]), .B(n28933), 
         .C(n33903), .D(n33904), .Z(n32196)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam \round_key_gen.trw_4__bdd_4_lut_28661 .init = 16'h6996;
    LUT4 i14536_3_lut_4_lut_4_lut (.A(n33846), .B(\round_logic.mixcolumns_block_71__N_1149[7] ), 
         .C(round_key[70]), .D(n33845), .Z(n13003)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14536_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 mux_692_Mux_60_i2_4_lut (.A(\round_key_gen.trw[4] ), .B(n7_adj_8139), 
         .C(n33846), .D(n8_adj_8137), .Z(n2_adj_8140)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_60_i2_4_lut.init = 16'h3aca;
    LUT4 \round_key_gen.trw_4__bdd_3_lut_28662  (.A(\round_key_gen.trw[4] ), 
         .B(n32196), .C(n33846), .Z(n32197)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \round_key_gen.trw_4__bdd_3_lut_28662 .init = 16'hcaca;
    PFUMX i28931 (.BLUT(n33217), .ALUT(n33216), .C0(n33847), .Z(n33218));
    LUT4 mux_692_Mux_61_i2_4_lut (.A(\round_key_gen.trw[5] ), .B(n7_adj_8141), 
         .C(n33846), .D(n8_adj_8142), .Z(n2_adj_8143)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_61_i2_4_lut.init = 16'h3aca;
    LUT4 mux_692_Mux_62_i2_4_lut (.A(\round_key_gen.trw[6] ), .B(n7_adj_8144), 
         .C(n33846), .D(n8_adj_8145), .Z(n2_adj_8146)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_62_i2_4_lut.init = 16'h3aca;
    LUT4 round_key_122__bdd_3_lut (.A(round_key[122]), .B(n33846), .C(\block_reg[0][26] ), 
         .Z(n32203)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_122__bdd_3_lut.init = 16'h4848;
    LUT4 \round_key_gen.trw_2__bdd_4_lut_28284  (.A(round_key[122]), .B(n33900), 
         .C(n33901), .D(\enc_new_block[82] ), .Z(n32205)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam \round_key_gen.trw_2__bdd_4_lut_28284 .init = 16'h6996;
    LUT4 \round_key_gen.trw_2__bdd_3_lut_28285  (.A(\round_key_gen.trw[2] ), 
         .B(n32205), .C(n33846), .Z(n32206)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \round_key_gen.trw_2__bdd_3_lut_28285 .init = 16'hcaca;
    LUT4 i14535_3_lut_4_lut_4_lut (.A(n33846), .B(\round_logic.mixcolumns_block_71__N_1149[0] ), 
         .C(round_key[71]), .D(n33845), .Z(n13004)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14535_3_lut_4_lut_4_lut.init = 16'h1400;
    FD1P3AX block_w1_reg__i1 (.D(n5291[64]), .SP(block_w1_we), .CK(clk_c), 
            .Q(\enc_new_block[64] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w1_reg__i1.GSR = "ENABLED";
    LUT4 mux_692_Mux_64_i2_4_lut (.A(\round_key_gen.trw[8] ), .B(n7_adj_8147), 
         .C(n33846), .D(n8_adj_8148), .Z(n2_adj_8149)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_64_i2_4_lut.init = 16'h3aca;
    PFUMX i28921 (.BLUT(n33205), .ALUT(n33204), .C0(n33847), .Z(n33206));
    LUT4 i14533_3_lut_4_lut_4_lut (.A(n33846), .B(\round_logic.mixcolumns_block_79__N_1341[2] ), 
         .C(round_key[73]), .D(n33845), .Z(n13006)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14533_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i14531_3_lut_4_lut_4_lut (.A(n33846), .B(\enc_new_block[11] ), 
         .C(round_key[75]), .D(n33845), .Z(n13008)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14531_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 mux_692_Mux_65_i2_4_lut (.A(\round_key_gen.trw[9] ), .B(n7_adj_8150), 
         .C(n33846), .D(n8_adj_8151), .Z(n2_adj_8152)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_65_i2_4_lut.init = 16'h3aca;
    LUT4 i14530_3_lut_4_lut_4_lut (.A(n33846), .B(\round_logic.mixcolumns_block_79__N_1341[5] ), 
         .C(round_key[76]), .D(n33845), .Z(n13009)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14530_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i14525_3_lut_4_lut_4_lut (.A(n33846), .B(\enc_new_block[49] ), 
         .C(round_key[81]), .D(n33845), .Z(n13014)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14525_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i14524_3_lut_4_lut_4_lut (.A(n33846), .B(\enc_new_block[50] ), 
         .C(round_key[82]), .D(n33845), .Z(n13015)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14524_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i14523_3_lut_4_lut_4_lut (.A(n33846), .B(\enc_new_block[51] ), 
         .C(round_key[83]), .D(n33845), .Z(n13016)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14523_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i14522_3_lut_4_lut_4_lut (.A(n33846), .B(\enc_new_block[52] ), 
         .C(round_key[84]), .D(n33845), .Z(n13017)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14522_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i14521_3_lut_4_lut_4_lut (.A(n33846), .B(\enc_new_block[53] ), 
         .C(round_key[85]), .D(n33845), .Z(n13018)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14521_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i14520_3_lut_4_lut_4_lut (.A(n33846), .B(\enc_new_block[54] ), 
         .C(round_key[86]), .D(n33845), .Z(n13019)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14520_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i14519_3_lut_4_lut_4_lut (.A(n33846), .B(\enc_new_block[55] ), 
         .C(round_key[87]), .D(n33845), .Z(n13020)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14519_3_lut_4_lut_4_lut.init = 16'h1400;
    PFUMX i28911 (.BLUT(n33193), .ALUT(n33192), .C0(n33847), .Z(n33194));
    LUT4 i1_2_lut_rep_565 (.A(\enc_new_block[60] ), .B(\enc_new_block[20] ), 
         .Z(n33869)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_rep_565.init = 16'h6666;
    LUT4 i14517_3_lut_4_lut_4_lut (.A(n33846), .B(\enc_new_block[89] ), 
         .C(round_key[89]), .D(n33845), .Z(n13022)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14517_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i14515_3_lut_4_lut_4_lut (.A(n33846), .B(\enc_new_block[91] ), 
         .C(round_key[91]), .D(n33845), .Z(n13024)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14515_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i14514_3_lut_4_lut_4_lut (.A(n33846), .B(\enc_new_block[92] ), 
         .C(round_key[92]), .D(n33845), .Z(n13025)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14514_3_lut_4_lut_4_lut.init = 16'h1400;
    FD1P3AX block_w2_reg__i1 (.D(n33072), .SP(block_w2_we), .CK(clk_c), 
            .Q(\enc_new_block[32] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w2_reg__i1.GSR = "ENABLED";
    LUT4 i1_4_lut (.A(n6347[3]), .B(n33841), .C(n20690), .D(n33847), 
         .Z(block_w2_we)) /* synthesis lut_function=(!(A+!(B (C+(D))+!B !((D)+!C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(422[7] 479[14])
    defparam i1_4_lut.init = 16'h4450;
    LUT4 i15168_3_lut (.A(n33845), .B(n33846), .C(block_w2_we_N_1489), 
         .Z(n20690)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i15168_3_lut.init = 16'hdcdc;
    LUT4 i14509_3_lut_4_lut_4_lut (.A(n33846), .B(\round_logic.mixcolumns_block_103__N_1101[2] ), 
         .C(round_key[97]), .D(n33845), .Z(n13030)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14509_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i14508_3_lut_4_lut_4_lut (.A(n33846), .B(\enc_new_block[2] ), .C(round_key[98]), 
         .D(n33845), .Z(n13031)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14508_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i14507_3_lut_4_lut_4_lut (.A(n33846), .B(\enc_new_block[3] ), .C(round_key[99]), 
         .D(n33845), .Z(n13032)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14507_3_lut_4_lut_4_lut.init = 16'h1400;
    FD1P3AY sword_ctr_reg_FSM_i0_i0 (.D(n25323), .SP(sword_ctr_we), .CK(clk_c), 
            .Q(n6364_c[0]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam sword_ctr_reg_FSM_i0_i0.GSR = "ENABLED";
    LUT4 i14504_3_lut_4_lut_4_lut (.A(n33846), .B(\round_logic.mixcolumns_block_103__N_1101[7] ), 
         .C(round_key[102]), .D(n33845), .Z(n13035)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14504_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i14501_3_lut_4_lut_4_lut (.A(n33846), .B(\round_logic.mixcolumns_block_111__N_1285[2] ), 
         .C(round_key[105]), .D(n33845), .Z(n13038)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14501_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i14499_3_lut_4_lut_4_lut (.A(n33846), .B(\enc_new_block[43] ), 
         .C(round_key[107]), .D(n33845), .Z(n13040)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14499_3_lut_4_lut_4_lut.init = 16'h1400;
    PFUMX i28900 (.BLUT(n33181), .ALUT(n33180), .C0(n33847), .Z(n33182));
    LUT4 i3_3_lut_4_lut_adj_333 (.A(\enc_new_block[60] ), .B(\enc_new_block[20] ), 
         .C(round_key[61]), .D(\round_logic.mixcolumns_block_39__N_1197[6] ), 
         .Z(n8_adj_8142)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i3_3_lut_4_lut_adj_333.init = 16'h6996;
    LUT4 i14498_3_lut_4_lut_4_lut (.A(n33846), .B(\round_logic.mixcolumns_block_111__N_1285[5] ), 
         .C(round_key[108]), .D(n33845), .Z(n13041)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14498_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i14493_3_lut_4_lut_4_lut (.A(n33846), .B(\enc_new_block[81] ), 
         .C(round_key[113]), .D(n33845), .Z(n13046)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14493_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 round_key_120__bdd_3_lut (.A(round_key[120]), .B(n33846), .C(\block_reg[0][24] ), 
         .Z(n32212)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_120__bdd_3_lut.init = 16'h4848;
    LUT4 mux_692_Mux_67_i2_4_lut (.A(\round_key_gen.trw[11] ), .B(n9_adj_8153), 
         .C(n33846), .D(n10_adj_8154), .Z(n2_adj_8155)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_67_i2_4_lut.init = 16'h3aca;
    LUT4 \round_key_gen.trw_0__bdd_4_lut_28371  (.A(round_key[120]), .B(n33903), 
         .C(n29077), .D(\enc_new_block[0] ), .Z(n32214)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam \round_key_gen.trw_0__bdd_4_lut_28371 .init = 16'h6996;
    LUT4 mux_692_Mux_68_i2_4_lut (.A(\round_key_gen.trw[12] ), .B(n7_adj_8156), 
         .C(n33846), .D(n8_adj_8157), .Z(n2_adj_8158)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_68_i2_4_lut.init = 16'h3aca;
    LUT4 \round_key_gen.trw_0__bdd_3_lut_28372  (.A(\round_key_gen.trw[0] ), 
         .B(n32214), .C(n33846), .Z(n32215)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \round_key_gen.trw_0__bdd_3_lut_28372 .init = 16'hcaca;
    PFUMX i28892 (.BLUT(n33172), .ALUT(n33171), .C0(n33847), .Z(n33173));
    LUT4 i14492_3_lut_4_lut_4_lut (.A(n33846), .B(\enc_new_block[82] ), 
         .C(round_key[114]), .D(n33845), .Z(n13047)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14492_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i14491_3_lut_4_lut_4_lut (.A(n33846), .B(\enc_new_block[83] ), 
         .C(round_key[115]), .D(n33845), .Z(n13048)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14491_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 mux_692_Mux_69_i2_4_lut (.A(\round_key_gen.trw[13] ), .B(n7_adj_8159), 
         .C(n33846), .D(n8_adj_8160), .Z(n2_adj_8161)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_69_i2_4_lut.init = 16'h3aca;
    LUT4 mux_692_Mux_70_i2_4_lut (.A(\round_key_gen.trw[14] ), .B(n7_adj_8162), 
         .C(n33846), .D(n8_adj_8163), .Z(n2_adj_8164)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_70_i2_4_lut.init = 16'h3aca;
    LUT4 n32180_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n32178), .D(n32180), 
         .Z(n32181)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n32180_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n32186_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n32184), .D(n32186), 
         .Z(n32187)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n32186_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n32197_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n32195), .D(n32197), 
         .Z(n32198)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n32197_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_692_Mux_71_i2_4_lut (.A(\round_key_gen.trw[15] ), .B(n7_adj_8165), 
         .C(n33846), .D(n8_adj_8166), .Z(n2_adj_8167)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_71_i2_4_lut.init = 16'h3aca;
    LUT4 n32206_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n32204), .D(n32206), 
         .Z(n32207)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n32206_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n32215_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n32213), .D(n32215), 
         .Z(n32216)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n32215_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n32227_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n32225), .D(n32227), 
         .Z(n32228)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n32227_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n32247_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n32245), .D(n32247), 
         .Z(n32248)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n32247_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n32253_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n32251), .D(n32253), 
         .Z(n32254)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n32253_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_692_Mux_73_i2_4_lut (.A(\round_key_gen.trw[17] ), .B(n7_adj_8168), 
         .C(n33846), .D(n8_adj_8169), .Z(n2_adj_8170)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_73_i2_4_lut.init = 16'h3aca;
    LUT4 n32259_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n32257), .D(n32259), 
         .Z(n32260)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n32259_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n32265_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n32263), .D(n32265), 
         .Z(n32266)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n32265_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 round_key_117__bdd_3_lut (.A(round_key[117]), .B(n33846), .C(\block_reg[0][21] ), 
         .Z(n32224)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_117__bdd_3_lut.init = 16'h4848;
    LUT4 new_sboxw_21__bdd_4_lut_28487 (.A(round_key[117]), .B(n33902), 
         .C(n29303), .D(\enc_new_block[125] ), .Z(n32226)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam new_sboxw_21__bdd_4_lut_28487.init = 16'h6996;
    LUT4 new_sboxw_21__bdd_3_lut_28488 (.A(\new_sboxw[21] ), .B(n32226), 
         .C(n33846), .Z(n32227)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam new_sboxw_21__bdd_3_lut_28488.init = 16'hcaca;
    LUT4 n32279_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n32277), .D(n32279), 
         .Z(n32280)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n32279_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n32288_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n32286), .D(n32288), 
         .Z(n32289)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n32288_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n32294_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n32292), .D(n32294), 
         .Z(n32295)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n32294_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n32303_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n32301), .D(n32303), 
         .Z(n32304)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n32303_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n32309_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n32307), .D(n32309), 
         .Z(n32310)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n32309_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n32324_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n32322), .D(n32324), 
         .Z(n32325)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n32324_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n32330_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n32328), .D(n32330), 
         .Z(n32331)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n32330_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n32336_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n32334), .D(n32336), 
         .Z(n32337)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n32336_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n32342_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n32340), .D(n32342), 
         .Z(n32343)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n32342_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n32366_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n32364), .D(n32366), 
         .Z(n32367)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n32366_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n32512_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n32510), .D(n32512), 
         .Z(n32513)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n32512_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n32558_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n32556), .D(n32558), 
         .Z(n32559)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n32558_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n32564_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n32562), .D(n32564), 
         .Z(n32565)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n32564_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n32575_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n32573), .D(n32575), 
         .Z(n32576)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n32575_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n32581_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n32579), .D(n32581), 
         .Z(n32582)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n32581_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n32604_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n32602), .D(n32604), 
         .Z(n32605)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n32604_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 round_key_112__bdd_3_lut (.A(round_key[112]), .B(n33846), .C(\block_reg[0][16] ), 
         .Z(n32244)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_112__bdd_3_lut.init = 16'h4848;
    LUT4 new_sboxw_16__bdd_4_lut_28410 (.A(round_key[112]), .B(n33895), 
         .C(n33896), .D(\enc_new_block[40] ), .Z(n32246)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam new_sboxw_16__bdd_4_lut_28410.init = 16'h6996;
    LUT4 new_sboxw_16__bdd_3_lut_28411 (.A(\new_sboxw[16] ), .B(n32246), 
         .C(n33846), .Z(n32247)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam new_sboxw_16__bdd_3_lut_28411.init = 16'hcaca;
    LUT4 round_key_111__bdd_3_lut (.A(round_key[111]), .B(n33846), .C(\block_reg[0][15] ), 
         .Z(n32250)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_111__bdd_3_lut.init = 16'h4848;
    LUT4 \round_key_gen.trw_23__bdd_4_lut_28415  (.A(round_key[111]), .B(n29399), 
         .C(n33907), .D(\enc_new_block[127] ), .Z(n32252)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam \round_key_gen.trw_23__bdd_4_lut_28415 .init = 16'h6996;
    LUT4 \round_key_gen.trw_23__bdd_3_lut_28416  (.A(\round_key_gen.trw[23] ), 
         .B(n32252), .C(n33846), .Z(n32253)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \round_key_gen.trw_23__bdd_3_lut_28416 .init = 16'hcaca;
    LUT4 round_key_110__bdd_3_lut (.A(round_key[110]), .B(n33846), .C(\block_reg[0][14] ), 
         .Z(n32256)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_110__bdd_3_lut.init = 16'h4848;
    LUT4 \round_key_gen.trw_22__bdd_4_lut_28423  (.A(round_key[110]), .B(n29303), 
         .C(n29037), .D(\enc_new_block[86] ), .Z(n32258)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam \round_key_gen.trw_22__bdd_4_lut_28423 .init = 16'h6996;
    LUT4 \round_key_gen.trw_22__bdd_3_lut_28424  (.A(\round_key_gen.trw[22] ), 
         .B(n32258), .C(n33846), .Z(n32259)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \round_key_gen.trw_22__bdd_3_lut_28424 .init = 16'hcaca;
    LUT4 round_key_109__bdd_3_lut (.A(round_key[109]), .B(n33846), .C(\block_reg[0][13] ), 
         .Z(n32262)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_109__bdd_3_lut.init = 16'h4848;
    LUT4 \round_key_gen.trw_21__bdd_4_lut_28428  (.A(round_key[109]), .B(n33852), 
         .C(\round_logic.mixcolumns_block_111__N_1285[5] ), .D(\round_logic.mixcolumns_block_103__N_1101[6] ), 
         .Z(n32264)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam \round_key_gen.trw_21__bdd_4_lut_28428 .init = 16'h6996;
    LUT4 \round_key_gen.trw_21__bdd_3_lut_28429  (.A(\round_key_gen.trw[21] ), 
         .B(n32264), .C(n33846), .Z(n32265)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \round_key_gen.trw_21__bdd_3_lut_28429 .init = 16'hcaca;
    LUT4 round_key_106__bdd_3_lut (.A(round_key[106]), .B(n33846), .C(\block_reg[0][10] ), 
         .Z(n32276)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_106__bdd_3_lut.init = 16'h4848;
    LUT4 \round_key_gen.trw_18__bdd_4_lut_28458  (.A(round_key[106]), .B(n33891), 
         .C(n33892), .D(\round_logic.mixcolumns_block_111__N_1285[2] ), 
         .Z(n32278)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam \round_key_gen.trw_18__bdd_4_lut_28458 .init = 16'h6996;
    LUT4 \round_key_gen.trw_18__bdd_3_lut_28448  (.A(\round_key_gen.trw[18] ), 
         .B(n32278), .C(n33846), .Z(n32279)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \round_key_gen.trw_18__bdd_3_lut_28448 .init = 16'hcaca;
    LUT4 round_key_104__bdd_3_lut_28450 (.A(round_key[104]), .B(n33846), 
         .C(\block_reg[0][8] ), .Z(n32285)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_104__bdd_3_lut_28450.init = 16'h4848;
    LUT4 \round_key_gen.trw_16__bdd_3_lut_28455  (.A(\round_key_gen.trw[16] ), 
         .B(n32287), .C(n33846), .Z(n32288)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \round_key_gen.trw_16__bdd_3_lut_28455 .init = 16'hcaca;
    LUT4 round_key_103__bdd_3_lut (.A(round_key[103]), .B(n33846), .C(\block_reg[0][7] ), 
         .Z(n32291)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_103__bdd_3_lut.init = 16'h4848;
    LUT4 n32701_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n32699), .D(n32701), 
         .Z(n32702)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n32701_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_692_Mux_75_i2_4_lut (.A(\round_key_gen.trw[19] ), .B(n7_adj_8171), 
         .C(n33846), .D(n8_adj_8172), .Z(n2_adj_8173)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_75_i2_4_lut.init = 16'h3aca;
    LUT4 mux_692_Mux_76_i2_4_lut (.A(\round_key_gen.trw[20] ), .B(n7_adj_8174), 
         .C(n33846), .D(n8_adj_8175), .Z(n2_adj_8176)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_76_i2_4_lut.init = 16'h3aca;
    LUT4 i4067_3_lut (.A(\enc_new_block[63] ), .B(\enc_new_block[31] ), 
         .C(n6364[3]), .Z(n9676)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam i4067_3_lut.init = 16'hcaca;
    LUT4 mux_178_i32_3_lut (.A(\enc_new_block[127] ), .B(\enc_new_block[95] ), 
         .C(n6364_c[1]), .Z(n2531[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam mux_178_i32_3_lut.init = 16'hcaca;
    LUT4 n32788_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n32786), .D(n32788), 
         .Z(n32789)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n32788_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n32854_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n32852), .D(n32854), 
         .Z(n32855)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n32854_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n32900_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n32898), .D(n32900), 
         .Z(n32901)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n32900_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i4065_3_lut (.A(\enc_new_block[62] ), .B(\enc_new_block[30] ), 
         .C(n6364[3]), .Z(n9674)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam i4065_3_lut.init = 16'hcaca;
    LUT4 n32913_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n32911), .D(n32913), 
         .Z(n32914)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n32913_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n32923_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n32921), .D(n32923), 
         .Z(n32924)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n32923_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n32937_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n32935), .D(n32937), 
         .Z(n32938)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n32937_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_178_i31_3_lut (.A(\enc_new_block[126] ), .B(\enc_new_block[94] ), 
         .C(n6364_c[1]), .Z(n2531[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam mux_178_i31_3_lut.init = 16'hcaca;
    LUT4 \round_key_gen.trw_15__bdd_4_lut_28378  (.A(round_key[103]), .B(n33896), 
         .C(n29037), .D(\enc_new_block[127] ), .Z(n32293)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam \round_key_gen.trw_15__bdd_4_lut_28378 .init = 16'h6996;
    LUT4 mux_692_Mux_81_i2_4_lut (.A(\new_sboxw[17] ), .B(n7_adj_8177), 
         .C(n33846), .D(n8_adj_8178), .Z(n2_adj_8179)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_81_i2_4_lut.init = 16'h3aca;
    LUT4 i4063_3_lut (.A(\enc_new_block[61] ), .B(\enc_new_block[29] ), 
         .C(n6364[3]), .Z(n9672)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam i4063_3_lut.init = 16'hcaca;
    LUT4 n32943_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n32941), .D(n32943), 
         .Z(n32944)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n32943_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n32952_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n32950), .D(n32952), 
         .Z(n32953)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n32952_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n32973_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n32971), .D(n32973), 
         .Z(n32974)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n32973_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_178_i30_3_lut (.A(\enc_new_block[125] ), .B(\enc_new_block[93] ), 
         .C(n6364_c[1]), .Z(n2531[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam mux_178_i30_3_lut.init = 16'hcaca;
    LUT4 n32982_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n32980), .D(n32982), 
         .Z(n32983)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n32982_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_692_Mux_82_i2_4_lut (.A(\new_sboxw[18] ), .B(n7_adj_8180), 
         .C(n33846), .D(n8_adj_8181), .Z(n2_adj_8182)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_82_i2_4_lut.init = 16'h3aca;
    LUT4 i4061_3_lut (.A(\enc_new_block[60] ), .B(\enc_new_block[28] ), 
         .C(n6364[3]), .Z(n9670)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam i4061_3_lut.init = 16'hcaca;
    LUT4 mux_178_i29_3_lut (.A(\enc_new_block[124] ), .B(\enc_new_block[92] ), 
         .C(n6364_c[1]), .Z(n2531[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam mux_178_i29_3_lut.init = 16'hcaca;
    LUT4 mux_692_Mux_83_i2_4_lut (.A(\new_sboxw[19] ), .B(n7_adj_8183), 
         .C(n33846), .D(n8_adj_8184), .Z(n2_adj_8185)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_83_i2_4_lut.init = 16'h3aca;
    LUT4 i4059_3_lut (.A(\enc_new_block[59] ), .B(\enc_new_block[27] ), 
         .C(n6364[3]), .Z(n9668)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam i4059_3_lut.init = 16'hcaca;
    LUT4 n32988_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n32986), .D(n32988), 
         .Z(n32989)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n32988_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_178_i28_3_lut (.A(\enc_new_block[123] ), .B(\enc_new_block[91] ), 
         .C(n6364_c[1]), .Z(n2531[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam mux_178_i28_3_lut.init = 16'hcaca;
    LUT4 n32997_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n32995), .D(n32997), 
         .Z(n32998)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n32997_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_692_Mux_84_i2_4_lut (.A(\new_sboxw[20] ), .B(n7_adj_8186), 
         .C(n33846), .D(n8_adj_8187), .Z(n2_adj_8188)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_84_i2_4_lut.init = 16'h3aca;
    LUT4 n33014_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n33012), .D(n33014), 
         .Z(n33015)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n33014_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i4057_3_lut (.A(\enc_new_block[58] ), .B(\enc_new_block[26] ), 
         .C(n6364[3]), .Z(n9666)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam i4057_3_lut.init = 16'hcaca;
    LUT4 n33026_bdd_3_lut_4_lut (.A(n33847), .B(n33845), .C(n33024), .D(n33026), 
         .Z(n33027)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam n33026_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 \round_key_gen.trw_15__bdd_3_lut_28379  (.A(\round_key_gen.trw[15] ), 
         .B(n32293), .C(n33846), .Z(n32294)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \round_key_gen.trw_15__bdd_3_lut_28379 .init = 16'hcaca;
    LUT4 mux_178_i27_3_lut (.A(\enc_new_block[122] ), .B(\enc_new_block[90] ), 
         .C(n6364_c[1]), .Z(n2531[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam mux_178_i27_3_lut.init = 16'hcaca;
    LUT4 mux_692_Mux_85_i2_4_lut (.A(\new_sboxw[21] ), .B(n7_adj_8189), 
         .C(n33846), .D(n8_adj_8190), .Z(n2_adj_8191)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_85_i2_4_lut.init = 16'h3aca;
    LUT4 i4055_3_lut (.A(\enc_new_block[57] ), .B(\enc_new_block[25] ), 
         .C(n6364[3]), .Z(n9664)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam i4055_3_lut.init = 16'hcaca;
    LUT4 mux_692_Mux_86_i2_4_lut (.A(\new_sboxw[22] ), .B(n7_adj_8192), 
         .C(n33846), .D(n8_adj_8193), .Z(n2_adj_8194)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_86_i2_4_lut.init = 16'h3aca;
    LUT4 mux_178_i26_3_lut (.A(\enc_new_block[121] ), .B(\enc_new_block[89] ), 
         .C(n6364_c[1]), .Z(n2531[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam mux_178_i26_3_lut.init = 16'hcaca;
    LUT4 mux_692_Mux_87_i2_4_lut (.A(\new_sboxw[23] ), .B(n7_adj_8195), 
         .C(n33846), .D(n8_adj_8196), .Z(n2_adj_8197)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_87_i2_4_lut.init = 16'h3aca;
    PFUMX i28882 (.BLUT(n33158), .ALUT(n33157), .C0(n33847), .Z(n33159));
    LUT4 i1_2_lut_rep_566 (.A(\enc_new_block[21] ), .B(\round_logic.mixcolumns_block_47__N_1397[7] ), 
         .Z(n33870)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_rep_566.init = 16'h6666;
    LUT4 i14490_3_lut_4_lut_4_lut (.A(n33846), .B(\enc_new_block[84] ), 
         .C(round_key[116]), .D(n33845), .Z(n13049)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14490_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i14488_3_lut_4_lut_4_lut (.A(n33846), .B(\enc_new_block[86] ), 
         .C(round_key[118]), .D(n33845), .Z(n13051)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14488_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i14487_3_lut_4_lut_4_lut (.A(n33846), .B(\enc_new_block[87] ), 
         .C(round_key[119]), .D(n33845), .Z(n13052)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14487_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i14485_3_lut_4_lut_4_lut (.A(n33846), .B(\enc_new_block[121] ), 
         .C(round_key[121]), .D(n33845), .Z(n13054)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14485_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i14483_3_lut_4_lut_4_lut (.A(n33846), .B(\enc_new_block[123] ), 
         .C(round_key[123]), .D(n33845), .Z(n13056)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14483_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 round_key_126__bdd_3_lut_28156_4_lut_4_lut (.A(n33846), .B(round_key[126]), 
         .C(\enc_new_block[126] ), .D(n33845), .Z(n32182)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_126__bdd_3_lut_28156_4_lut_4_lut.init = 16'h1400;
    LUT4 round_key_124__bdd_3_lut_28163_4_lut_4_lut (.A(n33846), .B(round_key[124]), 
         .C(\enc_new_block[124] ), .D(n33845), .Z(n32193)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_124__bdd_3_lut_28163_4_lut_4_lut.init = 16'h1400;
    LUT4 round_key_127__bdd_3_lut_28153_4_lut_4_lut (.A(n33846), .B(round_key[127]), 
         .C(\enc_new_block[127] ), .D(n33845), .Z(n32176)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam round_key_127__bdd_3_lut_28153_4_lut_4_lut.init = 16'h1400;
    LUT4 i15416_3_lut_4_lut_4_lut (.A(n33846), .B(\round_logic.mixcolumns_block_7__N_1245[2] ), 
         .C(round_key[1]), .D(n33845), .Z(n12934)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i15416_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i15415_3_lut_4_lut_4_lut (.A(n33846), .B(\enc_new_block[34] ), 
         .C(round_key[2]), .D(n33845), .Z(n12935)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i15415_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i15414_3_lut_4_lut_4_lut (.A(n33846), .B(\enc_new_block[35] ), 
         .C(round_key[3]), .D(n33845), .Z(n12936)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i15414_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i15413_3_lut_4_lut_4_lut (.A(n33846), .B(\round_logic.mixcolumns_block_7__N_1245[5] ), 
         .C(round_key[4]), .D(n33845), .Z(n12937)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i15413_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i15411_3_lut_4_lut_4_lut (.A(n33846), .B(\round_logic.mixcolumns_block_7__N_1245[6] ), 
         .C(round_key[5]), .D(n33845), .Z(n12938)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i15411_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i15409_3_lut_4_lut_4_lut (.A(n33846), .B(\round_logic.mixcolumns_block_7__N_1245[0] ), 
         .C(round_key[7]), .D(n33845), .Z(n12940)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i15409_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i15406_3_lut_4_lut_4_lut (.A(n33846), .B(\enc_new_block[74] ), 
         .C(round_key[10]), .D(n33845), .Z(n12943)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i15406_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i15404_3_lut_4_lut_4_lut (.A(n33846), .B(\round_logic.mixcolumns_block_15__N_1453[5] ), 
         .C(round_key[12]), .D(n33845), .Z(n12945)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i15404_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i15402_3_lut_4_lut_4_lut (.A(n33846), .B(\round_logic.mixcolumns_block_15__N_1453[7] ), 
         .C(round_key[14]), .D(n33845), .Z(n12947)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i15402_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i15399_3_lut_4_lut_4_lut (.A(n33846), .B(\enc_new_block[113] ), 
         .C(round_key[17]), .D(n33845), .Z(n12950)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i15399_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i15397_3_lut_4_lut_4_lut (.A(n33846), .B(\enc_new_block[115] ), 
         .C(round_key[19]), .D(n33845), .Z(n12952)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i15397_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i15396_3_lut_4_lut_4_lut (.A(n33846), .B(\enc_new_block[116] ), 
         .C(round_key[20]), .D(n33845), .Z(n12953)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i15396_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i3_3_lut_4_lut_adj_334 (.A(\enc_new_block[21] ), .B(\round_logic.mixcolumns_block_47__N_1397[7] ), 
         .C(\enc_new_block[22] ), .D(\enc_new_block[61] ), .Z(n8_adj_8145)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i3_3_lut_4_lut_adj_334.init = 16'h6996;
    LUT4 i15395_3_lut_4_lut_4_lut (.A(n33846), .B(\enc_new_block[117] ), 
         .C(round_key[21]), .D(n33845), .Z(n12954)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i15395_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i15391_3_lut_4_lut_4_lut (.A(n33846), .B(\enc_new_block[25] ), 
         .C(round_key[25]), .D(n33845), .Z(n12958)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i15391_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i14481_3_lut_4_lut_4_lut (.A(n33846), .B(\enc_new_block[125] ), 
         .C(round_key[125]), .D(n33845), .Z(n13058)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(331[9:21])
    defparam i14481_3_lut_4_lut_4_lut.init = 16'h1400;
    LUT4 i1_2_lut_rep_567 (.A(\round_logic.mixcolumns_block_39__N_1197[0] ), 
         .B(\round_logic.mixcolumns_block_47__N_1397[0] ), .Z(n33871)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i1_2_lut_rep_567.init = 16'h6666;
    LUT4 \round_key_gen.trw_0__bdd_3_lut_28541  (.A(\round_key_gen.trw[0] ), 
         .B(n32511), .C(n33846), .Z(n32512)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \round_key_gen.trw_0__bdd_3_lut_28541 .init = 16'hcaca;
    PFUMX i28862 (.BLUT(n33137), .ALUT(n33136), .C0(n33847), .Z(n33138));
    PFUMX i28857 (.BLUT(n33131), .ALUT(n33130), .C0(n33847), .Z(n33132));
    LUT4 i1_2_lut_rep_568 (.A(\enc_new_block[88] ), .B(\enc_new_block[96] ), 
         .Z(n33872)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_rep_568.init = 16'h6666;
    PFUMX i28849 (.BLUT(n33122), .ALUT(n33121), .C0(n33847), .Z(n33123));
    PFUMX i28837 (.BLUT(n33108), .ALUT(n33107), .C0(n33847), .Z(n33109));
    LUT4 \round_key_gen.trw_0__bdd_4_lut_28540  (.A(round_key[88]), .B(n33882), 
         .C(n29058), .D(\enc_new_block[48] ), .Z(n32511)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam \round_key_gen.trw_0__bdd_4_lut_28540 .init = 16'h6996;
    LUT4 i27501_3_lut_4_lut (.A(\block_new_127__N_1645[125] ), .B(n33846), 
         .C(n33847), .D(n13058), .Z(n5932[125])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27501_3_lut_4_lut.init = 16'hf808;
    LUT4 i27497_3_lut_4_lut (.A(\block_new_127__N_1645[123] ), .B(n33846), 
         .C(n33847), .D(n13056), .Z(n5932[123])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27497_3_lut_4_lut.init = 16'hf808;
    LUT4 i27493_3_lut_4_lut (.A(\block_new_127__N_1645[121] ), .B(n33846), 
         .C(n33847), .D(n13054), .Z(n5932[121])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27493_3_lut_4_lut.init = 16'hf808;
    LUT4 i27489_3_lut_4_lut (.A(\block_new_127__N_1645[119] ), .B(n33846), 
         .C(n33847), .D(n13052), .Z(n5932[119])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27489_3_lut_4_lut.init = 16'hf808;
    LUT4 round_key_88__bdd_3_lut (.A(round_key[88]), .B(n33846), .C(\block_reg[1][24] ), 
         .Z(n32509)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_88__bdd_3_lut.init = 16'h4848;
    LUT4 i27487_3_lut_4_lut (.A(\block_new_127__N_1645[118] ), .B(n33846), 
         .C(n33847), .D(n13051), .Z(n5932[118])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27487_3_lut_4_lut.init = 16'hf808;
    LUT4 i27483_3_lut_4_lut (.A(\block_new_127__N_1645[116] ), .B(n33846), 
         .C(n33847), .D(n13049), .Z(n5932[116])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27483_3_lut_4_lut.init = 16'hf808;
    LUT4 i27481_3_lut_4_lut (.A(\block_new_127__N_1645[115] ), .B(n33846), 
         .C(n33847), .D(n13048), .Z(n5932[115])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27481_3_lut_4_lut.init = 16'hf808;
    PFUMX i28821 (.BLUT(n33089), .ALUT(n33088), .C0(n33847), .Z(n33090));
    LUT4 i27479_3_lut_4_lut (.A(\block_new_127__N_1645[114] ), .B(n33846), 
         .C(n33847), .D(n13047), .Z(n5932[114])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27479_3_lut_4_lut.init = 16'hf808;
    LUT4 i27477_3_lut_4_lut (.A(\block_new_127__N_1645[113] ), .B(n33846), 
         .C(n33847), .D(n13046), .Z(n5932[113])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27477_3_lut_4_lut.init = 16'hf808;
    PFUMX i28812 (.BLUT(n33077), .ALUT(n33076), .C0(n33847), .Z(n33078));
    LUT4 i27467_3_lut_4_lut (.A(\block_new_127__N_1645[108] ), .B(n33846), 
         .C(n33847), .D(n13041), .Z(n5932[108])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27467_3_lut_4_lut.init = 16'hf808;
    LUT4 round_key_80__bdd_3_lut (.A(round_key[80]), .B(n33846), .C(\block_reg[1][16] ), 
         .Z(n32555)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_80__bdd_3_lut.init = 16'h4848;
    LUT4 new_sboxw_16__bdd_4_lut_28474 (.A(round_key[80]), .B(n29058), .C(n33889), 
         .D(\enc_new_block[88] ), .Z(n32557)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam new_sboxw_16__bdd_4_lut_28474.init = 16'h6996;
    LUT4 new_sboxw_16__bdd_3_lut_28475 (.A(\new_sboxw[16] ), .B(n32557), 
         .C(n33846), .Z(n32558)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam new_sboxw_16__bdd_3_lut_28475.init = 16'hcaca;
    LUT4 round_key_79__bdd_3_lut (.A(round_key[79]), .B(n33846), .C(\block_reg[1][15] ), 
         .Z(n32561)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_79__bdd_3_lut.init = 16'h4848;
    LUT4 i27847_2_lut_rep_537_2_lut_4_lut (.A(n6347[1]), .B(n28866), .C(n33848), 
         .D(n33846), .Z(n33841)) /* synthesis lut_function=(!(A ((D)+!B)+!A (B (D)+!B ((D)+!C)))) */ ;
    defparam i27847_2_lut_rep_537_2_lut_4_lut.init = 16'h00dc;
    LUT4 \round_key_gen.trw_23__bdd_4_lut_28470  (.A(round_key[79]), .B(n33882), 
         .C(n33888), .D(\round_logic.mixcolumns_block_71__N_1149[0] ), .Z(n32563)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam \round_key_gen.trw_23__bdd_4_lut_28470 .init = 16'h6996;
    LUT4 \round_key_gen.trw_23__bdd_3_lut_28471  (.A(\round_key_gen.trw[23] ), 
         .B(n32563), .C(n33846), .Z(n32564)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \round_key_gen.trw_23__bdd_3_lut_28471 .init = 16'hcaca;
    LUT4 round_key_78__bdd_3_lut (.A(round_key[78]), .B(n33846), .C(\block_reg[1][14] ), 
         .Z(n32572)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_78__bdd_3_lut.init = 16'h4848;
    LUT4 \round_key_gen.trw_22__bdd_4_lut_28466  (.A(round_key[78]), .B(n33890), 
         .C(n33886), .D(\round_logic.mixcolumns_block_71__N_1149[7] ), .Z(n32574)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam \round_key_gen.trw_22__bdd_4_lut_28466 .init = 16'h6996;
    LUT4 \round_key_gen.trw_22__bdd_3_lut_28467  (.A(\round_key_gen.trw[22] ), 
         .B(n32574), .C(n33846), .Z(n32575)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \round_key_gen.trw_22__bdd_3_lut_28467 .init = 16'hcaca;
    LUT4 round_key_77__bdd_3_lut (.A(round_key[77]), .B(n33846), .C(\block_reg[1][13] ), 
         .Z(n32578)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_77__bdd_3_lut.init = 16'h4848;
    LUT4 \round_key_gen.trw_21__bdd_4_lut_28462  (.A(round_key[77]), .B(n33883), 
         .C(n33887), .D(\round_logic.mixcolumns_block_71__N_1149[6] ), .Z(n32580)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam \round_key_gen.trw_21__bdd_4_lut_28462 .init = 16'h6996;
    LUT4 \round_key_gen.trw_21__bdd_3_lut_28463  (.A(\round_key_gen.trw[21] ), 
         .B(n32580), .C(n33846), .Z(n32581)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \round_key_gen.trw_21__bdd_3_lut_28463 .init = 16'hcaca;
    LUT4 i27465_3_lut_4_lut (.A(\block_new_127__N_1645[107] ), .B(n33846), 
         .C(n33847), .D(n13040), .Z(n5932[107])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27465_3_lut_4_lut.init = 16'hf808;
    LUT4 i27461_3_lut_4_lut (.A(\block_new_127__N_1645[105] ), .B(n33846), 
         .C(n33847), .D(n13038), .Z(n5932[105])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27461_3_lut_4_lut.init = 16'hf808;
    LUT4 i27455_3_lut_4_lut (.A(\block_new_127__N_1645[102] ), .B(n33846), 
         .C(n33847), .D(n13035), .Z(n5932[102])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27455_3_lut_4_lut.init = 16'hf808;
    LUT4 round_key_74__bdd_3_lut (.A(round_key[74]), .B(n33846), .C(\block_reg[1][10] ), 
         .Z(n32601)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_74__bdd_3_lut.init = 16'h4848;
    LUT4 \round_key_gen.trw_18__bdd_3_lut_28459  (.A(\round_key_gen.trw[18] ), 
         .B(n32603), .C(n33846), .Z(n32604)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \round_key_gen.trw_18__bdd_3_lut_28459 .init = 16'hcaca;
    LUT4 i27449_3_lut_4_lut (.A(\block_new_127__N_1645[99] ), .B(n33846), 
         .C(n33847), .D(n13032), .Z(n5932[99])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27449_3_lut_4_lut.init = 16'hf808;
    LUT4 i3_3_lut_4_lut_adj_335 (.A(\enc_new_block[88] ), .B(\enc_new_block[96] ), 
         .C(\round_logic.mixcolumns_block_79__N_1341[2] ), .D(round_key[65]), 
         .Z(n8_adj_8151)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i3_3_lut_4_lut_adj_335.init = 16'h6996;
    PFUMX i28806 (.BLUT(n33068), .ALUT(n33067), .C0(n33847), .Z(n33069));
    LUT4 i27447_3_lut_4_lut (.A(\block_new_127__N_1645[98] ), .B(n33846), 
         .C(n33847), .D(n13031), .Z(n5932[98])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27447_3_lut_4_lut.init = 16'hf808;
    LUT4 i27445_3_lut_4_lut (.A(\block_new_127__N_1645[97] ), .B(n33846), 
         .C(n33847), .D(n13030), .Z(n5932[97])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27445_3_lut_4_lut.init = 16'hf808;
    LUT4 round_key_72__bdd_3_lut (.A(round_key[72]), .B(n33846), .C(\block_reg[1][8] ), 
         .Z(n32698)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_72__bdd_3_lut.init = 16'h4848;
    LUT4 \round_key_gen.trw_16__bdd_4_lut_29731  (.A(round_key[72]), .B(n33875), 
         .C(n33872), .D(\enc_new_block[48] ), .Z(n32700)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam \round_key_gen.trw_16__bdd_4_lut_29731 .init = 16'h6996;
    LUT4 \round_key_gen.trw_16__bdd_3_lut_28769  (.A(\round_key_gen.trw[16] ), 
         .B(n32700), .C(n33846), .Z(n32701)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \round_key_gen.trw_16__bdd_3_lut_28769 .init = 16'hcaca;
    LUT4 round_key_35__bdd_3_lut (.A(round_key[35]), .B(n33846), .C(\block_reg[2][3] ), 
         .Z(n33053)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_35__bdd_3_lut.init = 16'h4848;
    LUT4 \round_key_gen.trw_11__bdd_3_lut  (.A(\round_key_gen.trw[11] ), .B(n33055), 
         .C(n33846), .Z(n33056)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \round_key_gen.trw_11__bdd_3_lut .init = 16'hcaca;
    LUT4 i1_2_lut_rep_571 (.A(\round_logic.mixcolumns_block_71__N_1149[0] ), 
         .B(\round_logic.mixcolumns_block_79__N_1341[0] ), .Z(n33875)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i1_2_lut_rep_571.init = 16'h6666;
    LUT4 i1_3_lut_rep_541_4_lut (.A(enc_round_nr[3]), .B(n33914), .C(n28866), 
         .D(n6347[1]), .Z(n33845)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A (C)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(387[27:47])
    defparam i1_3_lut_rep_541_4_lut.init = 16'hf0f8;
    LUT4 i1_3_lut_4_lut (.A(enc_round_nr[3]), .B(n33914), .C(n6347[2]), 
         .D(n6347[0]), .Z(n2924)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A (C+(D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(387[27:47])
    defparam i1_3_lut_4_lut.init = 16'hf7f0;
    LUT4 i27874_3_lut_rep_543_4_lut (.A(enc_round_nr[3]), .B(n33914), .C(n6347[1]), 
         .D(n28866), .Z(n33847)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(387[27:47])
    defparam i27874_3_lut_rep_543_4_lut.init = 16'h0008;
    LUT4 i27891_2_lut_rep_539_4_lut_3_lut_4_lut (.A(enc_round_nr[3]), .B(n33914), 
         .C(n6347[1]), .D(n28866), .Z(n33843)) /* synthesis lut_function=(A (B ((D)+!C)+!B (D))+!A (D)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(387[27:47])
    defparam i27891_2_lut_rep_539_4_lut_3_lut_4_lut.init = 16'hff08;
    LUT4 i27435_3_lut_4_lut (.A(\block_new_127__N_1645[92] ), .B(n33846), 
         .C(n33847), .D(n13025), .Z(n5932[92])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27435_3_lut_4_lut.init = 16'hf808;
    LUT4 i27433_3_lut_4_lut (.A(\block_new_127__N_1645[91] ), .B(n33846), 
         .C(n33847), .D(n13024), .Z(n5932[91])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27433_3_lut_4_lut.init = 16'hf808;
    LUT4 i27429_3_lut_4_lut (.A(\block_new_127__N_1645[89] ), .B(n33846), 
         .C(n33847), .D(n13022), .Z(n5932[89])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27429_3_lut_4_lut.init = 16'hf808;
    LUT4 i27425_3_lut_4_lut (.A(\block_new_127__N_1645[87] ), .B(n33846), 
         .C(n33847), .D(n13020), .Z(n5932[87])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27425_3_lut_4_lut.init = 16'hf808;
    LUT4 i27423_3_lut_4_lut (.A(\block_new_127__N_1645[86] ), .B(n33846), 
         .C(n33847), .D(n13019), .Z(n5932[86])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27423_3_lut_4_lut.init = 16'hf808;
    LUT4 i27421_3_lut_4_lut (.A(\block_new_127__N_1645[85] ), .B(n33846), 
         .C(n33847), .D(n13018), .Z(n5932[85])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27421_3_lut_4_lut.init = 16'hf808;
    LUT4 i27419_3_lut_4_lut (.A(\block_new_127__N_1645[84] ), .B(n33846), 
         .C(n33847), .D(n13017), .Z(n5932[84])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27419_3_lut_4_lut.init = 16'hf808;
    LUT4 round_key_66__bdd_3_lut (.A(round_key[66]), .B(n33846), .C(\block_reg[1][2] ), 
         .Z(n32785)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_66__bdd_3_lut.init = 16'h4848;
    LUT4 i27417_3_lut_4_lut (.A(\block_new_127__N_1645[83] ), .B(n33846), 
         .C(n33847), .D(n13016), .Z(n5932[83])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27417_3_lut_4_lut.init = 16'hf808;
    LUT4 i27415_3_lut_4_lut (.A(\block_new_127__N_1645[82] ), .B(n33846), 
         .C(n33847), .D(n13015), .Z(n5932[82])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27415_3_lut_4_lut.init = 16'hf808;
    LUT4 i3_3_lut_4_lut_adj_336 (.A(\round_logic.mixcolumns_block_71__N_1149[0] ), 
         .B(\round_logic.mixcolumns_block_79__N_1341[0] ), .C(round_key[76]), 
         .D(n33881), .Z(n8_adj_8175)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i3_3_lut_4_lut_adj_336.init = 16'h6996;
    LUT4 i3_3_lut_4_lut_adj_337 (.A(\round_logic.mixcolumns_block_71__N_1149[0] ), 
         .B(\round_logic.mixcolumns_block_79__N_1341[0] ), .C(\round_logic.mixcolumns_block_71__N_1149[2] ), 
         .D(n29058), .Z(n8_adj_8169)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i3_3_lut_4_lut_adj_337.init = 16'h6996;
    LUT4 i1_2_lut_rep_572 (.A(\round_logic.mixcolumns_block_79__N_1341[2] ), 
         .B(\enc_new_block[98] ), .Z(n33876)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_rep_572.init = 16'h6666;
    LUT4 i3_3_lut_4_lut_adj_338 (.A(\round_logic.mixcolumns_block_79__N_1341[2] ), 
         .B(\enc_new_block[98] ), .C(\enc_new_block[49] ), .D(\enc_new_block[90] ), 
         .Z(n8_adj_8181)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i3_3_lut_4_lut_adj_338.init = 16'h6996;
    LUT4 i2_2_lut (.A(\enc_new_block[17] ), .B(\enc_new_block[58] ), .Z(n7_adj_8128)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i2_2_lut.init = 16'h6666;
    LUT4 \round_key_gen.trw_10__bdd_4_lut_29765  (.A(round_key[66]), .B(n33851), 
         .C(\enc_new_block[89] ), .D(\enc_new_block[10] ), .Z(n32787)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam \round_key_gen.trw_10__bdd_4_lut_29765 .init = 16'h6996;
    LUT4 \round_key_gen.trw_10__bdd_3_lut  (.A(\round_key_gen.trw[10] ), .B(n32787), 
         .C(n33846), .Z(n32788)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \round_key_gen.trw_10__bdd_3_lut .init = 16'hcaca;
    LUT4 i1_2_lut (.A(\enc_new_block[64] ), .B(\enc_new_block[56] ), .Z(n29071)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut.init = 16'h6666;
    LUT4 i27413_3_lut_4_lut (.A(\block_new_127__N_1645[81] ), .B(n33846), 
         .C(n33847), .D(n13014), .Z(n5932[81])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27413_3_lut_4_lut.init = 16'hf808;
    LUT4 i2_2_lut_adj_339 (.A(\enc_new_block[107] ), .B(\round_logic.mixcolumns_block_39__N_1197[5] ), 
         .Z(n7_adj_8120)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i2_2_lut_adj_339.init = 16'h6666;
    LUT4 i2_2_lut_adj_340 (.A(\enc_new_block[19] ), .B(\enc_new_block[59] ), 
         .Z(n7_adj_8117)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i2_2_lut_adj_340.init = 16'h6666;
    LUT4 i2_2_lut_adj_341 (.A(round_key[41]), .B(\round_logic.mixcolumns_block_39__N_1197[2] ), 
         .Z(n7_adj_8105)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i2_2_lut_adj_341.init = 16'h6666;
    LUT4 i2_2_lut_adj_342 (.A(\enc_new_block[63] ), .B(\enc_new_block[62] ), 
         .Z(n7_adj_8096)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i2_2_lut_adj_342.init = 16'h6666;
    LUT4 i2_2_lut_adj_343 (.A(\enc_new_block[60] ), .B(round_key[37]), .Z(n7_adj_8081)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i2_2_lut_adj_343.init = 16'h6666;
    LUT4 i27403_3_lut_4_lut (.A(\block_new_127__N_1645[76] ), .B(n33846), 
         .C(n33847), .D(n13009), .Z(n5932[76])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27403_3_lut_4_lut.init = 16'hf808;
    LUT4 round_key_63__bdd_3_lut (.A(round_key[63]), .B(n33846), .C(\block_reg[2][31] ), 
         .Z(n32851)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_63__bdd_3_lut.init = 16'h4848;
    LUT4 i27401_3_lut_4_lut (.A(\block_new_127__N_1645[75] ), .B(n33846), 
         .C(n33847), .D(n13008), .Z(n5932[75])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27401_3_lut_4_lut.init = 16'hf808;
    LUT4 i27397_3_lut_4_lut (.A(\block_new_127__N_1645[73] ), .B(n33846), 
         .C(n33847), .D(n13006), .Z(n5932[73])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27397_3_lut_4_lut.init = 16'hf808;
    LUT4 i2_2_lut_adj_344 (.A(round_key[36]), .B(\round_logic.mixcolumns_block_47__N_1397[5] ), 
         .Z(n7_adj_8062)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i2_2_lut_adj_344.init = 16'h6666;
    LUT4 i4_4_lut (.A(n33862), .B(\enc_new_block[59] ), .C(\enc_new_block[58] ), 
         .D(\enc_new_block[66] ), .Z(n10_adj_8123)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i4_4_lut.init = 16'h6996;
    LUT4 i2_2_lut_adj_345 (.A(round_key[34]), .B(\enc_new_block[106] ), 
         .Z(n7_adj_8053)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i2_2_lut_adj_345.init = 16'h6666;
    LUT4 i2_2_lut_adj_346 (.A(round_key[33]), .B(\round_logic.mixcolumns_block_47__N_1397[2] ), 
         .Z(n7_adj_8050)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i2_2_lut_adj_346.init = 16'h6666;
    LUT4 i2_2_lut_adj_347 (.A(round_key[30]), .B(\enc_new_block[117] ), 
         .Z(n7_adj_8047)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i2_2_lut_adj_347.init = 16'h6666;
    LUT4 \round_key_gen.trw_7__bdd_4_lut_28699  (.A(round_key[63]), .B(n33871), 
         .C(n11620), .D(\enc_new_block[23] ), .Z(n32853)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam \round_key_gen.trw_7__bdd_4_lut_28699 .init = 16'h6996;
    LUT4 \round_key_gen.trw_18__bdd_3_lut_28449_4_lut  (.A(\round_logic.mixcolumns_block_71__N_1149[2] ), 
         .B(n33880), .C(n33876), .D(round_key[74]), .Z(n32603)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam \round_key_gen.trw_18__bdd_3_lut_28449_4_lut .init = 16'h6996;
    LUT4 i3_3_lut_4_lut_adj_348 (.A(\enc_new_block[11] ), .B(n33889), .C(n33883), 
         .D(\enc_new_block[51] ), .Z(n8_adj_8187)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i3_3_lut_4_lut_adj_348.init = 16'h6996;
    LUT4 i3_3_lut_4_lut_adj_349 (.A(\enc_new_block[11] ), .B(n33889), .C(round_key[83]), 
         .D(\enc_new_block[50] ), .Z(n8_adj_8184)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i3_3_lut_4_lut_adj_349.init = 16'h6996;
    LUT4 i3_3_lut_4_lut_adj_350 (.A(\enc_new_block[0] ), .B(n33894), .C(round_key[105]), 
         .D(\round_logic.mixcolumns_block_103__N_1101[2] ), .Z(n8_adj_8072)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i3_3_lut_4_lut_adj_350.init = 16'h6996;
    LUT4 \round_key_gen.trw_16__bdd_3_lut_28228_4_lut  (.A(\enc_new_block[0] ), 
         .B(n33894), .C(n33898), .D(round_key[104]), .Z(n32287)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam \round_key_gen.trw_16__bdd_3_lut_28228_4_lut .init = 16'h6996;
    LUT4 \round_key_gen.trw_7__bdd_3_lut_28700  (.A(\round_key_gen.trw[7] ), 
         .B(n32853), .C(n33846), .Z(n32854)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \round_key_gen.trw_7__bdd_3_lut_28700 .init = 16'hcaca;
    LUT4 \round_key_gen.trw_13__bdd_3_lut_28238_4_lut  (.A(\round_logic.mixcolumns_block_103__N_1101[5] ), 
         .B(n33906), .C(n33905), .D(round_key[101]), .Z(n32302)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam \round_key_gen.trw_13__bdd_3_lut_28238_4_lut .init = 16'h6996;
    LUT4 i1_2_lut_adj_351 (.A(\enc_new_block[28] ), .B(\enc_new_block[116] ), 
         .Z(n11634)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_adj_351.init = 16'h6666;
    LUT4 i27393_3_lut_4_lut (.A(\block_new_127__N_1645[71] ), .B(n33846), 
         .C(n33847), .D(n13004), .Z(n5932[71])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27393_3_lut_4_lut.init = 16'hf808;
    LUT4 i4_4_lut_adj_352 (.A(\enc_new_block[116] ), .B(round_key[28]), 
         .C(\enc_new_block[115] ), .D(\round_logic.mixcolumns_block_7__N_1245[5] ), 
         .Z(n10_adj_8045)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i4_4_lut_adj_352.init = 16'h6996;
    LUT4 i1_2_lut_adj_353 (.A(\enc_new_block[34] ), .B(\enc_new_block[74] ), 
         .Z(n11641)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_adj_353.init = 16'h6666;
    LUT4 i1_2_lut_adj_354 (.A(\enc_new_block[25] ), .B(\enc_new_block[113] ), 
         .Z(n11630)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_adj_354.init = 16'h6666;
    LUT4 i3_2_lut (.A(\enc_new_block[113] ), .B(\round_logic.mixcolumns_block_7__N_1245[2] ), 
         .Z(n9)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i3_2_lut.init = 16'h6666;
    LUT4 i4_4_lut_adj_355 (.A(n33926), .B(n12156), .C(\round_logic.mixcolumns_block_15__N_1453[2] ), 
         .D(round_key[25]), .Z(n10)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i4_4_lut_adj_355.init = 16'h6996;
    LUT4 i1_2_lut_adj_356 (.A(\enc_new_block[24] ), .B(\enc_new_block[112] ), 
         .Z(n12156)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_adj_356.init = 16'h6666;
    LUT4 i1_2_lut_adj_357 (.A(\enc_new_block[72] ), .B(\enc_new_block[32] ), 
         .Z(n29080)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_adj_357.init = 16'h6666;
    LUT4 i2_2_lut_adj_358 (.A(\enc_new_block[116] ), .B(\round_logic.mixcolumns_block_15__N_1453[5] ), 
         .Z(n7_adj_8028)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i2_2_lut_adj_358.init = 16'h6666;
    LUT4 i4_4_lut_adj_359 (.A(\round_logic.mixcolumns_block_15__N_1453[0] ), 
         .B(\enc_new_block[25] ), .C(\round_logic.mixcolumns_block_15__N_1453[2] ), 
         .D(round_key[17]), .Z(n10_adj_8198)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i4_4_lut_adj_359.init = 16'h6996;
    LUT4 i2_2_lut_adj_360 (.A(\round_logic.mixcolumns_block_7__N_1245[7] ), 
         .B(\round_logic.mixcolumns_block_15__N_1453[6] ), .Z(n7_adj_8199)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i2_2_lut_adj_360.init = 16'h6666;
    LUT4 i4_4_lut_adj_361 (.A(\enc_new_block[115] ), .B(n11641), .C(\enc_new_block[35] ), 
         .D(\enc_new_block[27] ), .Z(n10_adj_8200)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i4_4_lut_adj_361.init = 16'h6996;
    LUT4 i2_2_lut_adj_362 (.A(\round_logic.mixcolumns_block_7__N_1245[2] ), 
         .B(\enc_new_block[114] ), .Z(n7_adj_8201)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i2_2_lut_adj_362.init = 16'h6666;
    LUT4 i27391_3_lut_4_lut (.A(\block_new_127__N_1645[70] ), .B(n33846), 
         .C(n33847), .D(n13003), .Z(n5932[70])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27391_3_lut_4_lut.init = 16'hf808;
    LUT4 i2_2_lut_adj_363 (.A(\enc_new_block[31] ), .B(\enc_new_block[30] ), 
         .Z(n7_adj_8202)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i2_2_lut_adj_363.init = 16'h6666;
    LUT4 round_key_58__bdd_3_lut (.A(round_key[58]), .B(n33846), .C(\block_reg[2][26] ), 
         .Z(n32897)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_58__bdd_3_lut.init = 16'h4848;
    LUT4 i2_2_lut_adj_364 (.A(\enc_new_block[28] ), .B(round_key[5]), .Z(n7_adj_8203)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i2_2_lut_adj_364.init = 16'h6666;
    LUT4 i2_2_lut_3_lut_adj_365 (.A(\enc_new_block[99] ), .B(\enc_new_block[91] ), 
         .C(\enc_new_block[10] ), .Z(n7_adj_8183)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i2_2_lut_3_lut_adj_365.init = 16'h9696;
    LUT4 i3_3_lut_4_lut_adj_366 (.A(\enc_new_block[99] ), .B(\enc_new_block[91] ), 
         .C(\enc_new_block[51] ), .D(round_key[75]), .Z(n8_adj_8172)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i3_3_lut_4_lut_adj_366.init = 16'h6996;
    LUT4 i3_3_lut_4_lut_adj_367 (.A(\enc_new_block[99] ), .B(\enc_new_block[91] ), 
         .C(round_key[68]), .D(n33877), .Z(n8_adj_8157)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i3_3_lut_4_lut_adj_367.init = 16'h6996;
    LUT4 i1_2_lut_rep_573 (.A(\round_logic.mixcolumns_block_71__N_1149[0] ), 
         .B(\enc_new_block[95] ), .Z(n33877)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i1_2_lut_rep_573.init = 16'h6666;
    LUT4 i3_3_lut_4_lut_adj_368 (.A(\round_logic.mixcolumns_block_71__N_1149[0] ), 
         .B(\enc_new_block[95] ), .C(\enc_new_block[54] ), .D(\round_logic.mixcolumns_block_79__N_1341[7] ), 
         .Z(n8_adj_8196)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i3_3_lut_4_lut_adj_368.init = 16'h6996;
    LUT4 i3_3_lut_4_lut_adj_369 (.A(\round_logic.mixcolumns_block_71__N_1149[0] ), 
         .B(\enc_new_block[95] ), .C(\enc_new_block[48] ), .D(round_key[64]), 
         .Z(n8_adj_8148)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i3_3_lut_4_lut_adj_369.init = 16'h6996;
    LUT4 i1_2_lut_rep_574 (.A(\enc_new_block[49] ), .B(\enc_new_block[89] ), 
         .Z(n33878)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_rep_574.init = 16'h6666;
    LUT4 i2_2_lut_adj_370 (.A(round_key[4]), .B(\enc_new_block[35] ), .Z(n7_adj_8204)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i2_2_lut_adj_370.init = 16'h6666;
    PFUMX i28793 (.BLUT(n33053), .ALUT(n33052), .C0(n33847), .Z(n33054));
    LUT4 i2_2_lut_adj_371 (.A(round_key[3]), .B(\enc_new_block[27] ), .Z(n7_adj_8205)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i2_2_lut_adj_371.init = 16'h6666;
    LUT4 i2_2_lut_adj_372 (.A(\enc_new_block[25] ), .B(round_key[2]), .Z(n7_adj_8206)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i2_2_lut_adj_372.init = 16'h6666;
    LUT4 i3_2_lut_adj_373 (.A(\round_logic.mixcolumns_block_15__N_1453[2] ), 
         .B(\enc_new_block[24] ), .Z(n9_adj_8207)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i3_2_lut_adj_373.init = 16'h6666;
    LUT4 i4_4_lut_adj_374 (.A(n33922), .B(n11630), .C(\enc_new_block[32] ), 
         .D(round_key[1]), .Z(n10_adj_8208)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i4_4_lut_adj_374.init = 16'h6996;
    LUT4 i2_2_lut_3_lut_4_lut (.A(\enc_new_block[49] ), .B(\enc_new_block[89] ), 
         .C(\enc_new_block[95] ), .D(\round_logic.mixcolumns_block_71__N_1149[0] ), 
         .Z(n7_adj_8150)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i2_2_lut_3_lut_4_lut.init = 16'h6996;
    LUT4 i2_2_lut_3_lut_adj_375 (.A(\enc_new_block[49] ), .B(\enc_new_block[89] ), 
         .C(round_key[73]), .Z(n7_adj_8168)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i2_2_lut_3_lut_adj_375.init = 16'h9696;
    LUT4 i1_2_lut_rep_575 (.A(\enc_new_block[98] ), .B(\enc_new_block[10] ), 
         .Z(n33879)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_rep_575.init = 16'h6666;
    LUT4 i2_2_lut_3_lut_4_lut_adj_376 (.A(\enc_new_block[98] ), .B(\enc_new_block[10] ), 
         .C(\round_logic.mixcolumns_block_79__N_1341[0] ), .D(\round_logic.mixcolumns_block_71__N_1149[0] ), 
         .Z(n7_adj_8171)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i2_2_lut_3_lut_4_lut_adj_376.init = 16'h6996;
    LUT4 i1_2_lut_rep_576 (.A(\enc_new_block[50] ), .B(\enc_new_block[90] ), 
         .Z(n33880)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i1_2_lut_rep_576.init = 16'h6666;
    LUT4 i1_2_lut_rep_547_3_lut (.A(\enc_new_block[50] ), .B(\enc_new_block[90] ), 
         .C(\round_logic.mixcolumns_block_71__N_1149[2] ), .Z(n33851)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i1_2_lut_rep_547_3_lut.init = 16'h9696;
    LUT4 i1_2_lut_rep_577 (.A(\enc_new_block[99] ), .B(\enc_new_block[11] ), 
         .Z(n33881)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i1_2_lut_rep_577.init = 16'h6666;
    LUT4 i3_3_lut_4_lut_adj_377 (.A(\enc_new_block[99] ), .B(\enc_new_block[11] ), 
         .C(\enc_new_block[51] ), .D(round_key[91]), .Z(n8_adj_8036)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i3_3_lut_4_lut_adj_377.init = 16'h6996;
    LUT4 i1_2_lut_rep_578 (.A(\enc_new_block[55] ), .B(\enc_new_block[95] ), 
         .Z(n33882)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i1_2_lut_rep_578.init = 16'h6666;
    LUT4 i2_2_lut_3_lut_adj_378 (.A(\enc_new_block[55] ), .B(\enc_new_block[95] ), 
         .C(\enc_new_block[52] ), .Z(n7_adj_8038)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i2_2_lut_3_lut_adj_378.init = 16'h9696;
    LUT4 i3_3_lut_4_lut_adj_379 (.A(\enc_new_block[55] ), .B(\enc_new_block[95] ), 
         .C(\enc_new_block[49] ), .D(n29083), .Z(n8_adj_8033)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i3_3_lut_4_lut_adj_379.init = 16'h6996;
    LUT4 i2_2_lut_3_lut_4_lut_adj_380 (.A(\enc_new_block[55] ), .B(\enc_new_block[95] ), 
         .C(\enc_new_block[90] ), .D(\enc_new_block[50] ), .Z(n7_adj_8035)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i2_2_lut_3_lut_4_lut_adj_380.init = 16'h6996;
    LUT4 i1_2_lut_rep_579 (.A(\round_logic.mixcolumns_block_79__N_1341[5] ), 
         .B(\round_logic.mixcolumns_block_71__N_1149[5] ), .Z(n33883)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_rep_579.init = 16'h6666;
    LUT4 i3_3_lut_4_lut_adj_381 (.A(\round_logic.mixcolumns_block_79__N_1341[5] ), 
         .B(\round_logic.mixcolumns_block_71__N_1149[5] ), .C(round_key[92]), 
         .D(n33884), .Z(n8_adj_8039)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i3_3_lut_4_lut_adj_381.init = 16'h6996;
    LUT4 i1_2_lut_rep_580 (.A(\enc_new_block[91] ), .B(\enc_new_block[51] ), 
         .Z(n33884)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i1_2_lut_rep_580.init = 16'h6666;
    LUT4 i3_2_lut_3_lut (.A(\enc_new_block[91] ), .B(\enc_new_block[51] ), 
         .C(\enc_new_block[98] ), .Z(n9_adj_8153)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i3_2_lut_3_lut.init = 16'h9696;
    LUT4 i1_2_lut_rep_581 (.A(\enc_new_block[52] ), .B(\enc_new_block[92] ), 
         .Z(n33885)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_rep_581.init = 16'h6666;
    LUT4 i2_2_lut_3_lut_adj_382 (.A(\enc_new_block[52] ), .B(\enc_new_block[92] ), 
         .C(\round_logic.mixcolumns_block_71__N_1149[5] ), .Z(n7_adj_8174)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i2_2_lut_3_lut_adj_382.init = 16'h9696;
    FD1P3AX enc_ctrl_reg_FSM_i0_i1 (.D(n2924), .SP(enc_ctrl_we), .CK(clk_c), 
            .Q(n6347[1]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(422[7] 479[14])
    defparam enc_ctrl_reg_FSM_i0_i1.GSR = "ENABLED";
    FD1P3AX enc_ctrl_reg_FSM_i0_i2 (.D(n33913), .SP(enc_ctrl_we), .CK(clk_c), 
            .Q(n6347[2]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(422[7] 479[14])
    defparam enc_ctrl_reg_FSM_i0_i2.GSR = "ENABLED";
    FD1P3AY enc_ctrl_reg_FSM_i0_i3 (.D(n28773), .SP(enc_ctrl_we), .CK(clk_c), 
            .Q(n6347[3]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(422[7] 479[14])
    defparam enc_ctrl_reg_FSM_i0_i3.GSR = "ENABLED";
    LUT4 i2_2_lut_3_lut_adj_383 (.A(\enc_new_block[52] ), .B(\enc_new_block[92] ), 
         .C(\round_logic.mixcolumns_block_79__N_1341[5] ), .Z(n7_adj_8156)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i2_2_lut_3_lut_adj_383.init = 16'h9696;
    LUT4 i1_2_lut_rep_582 (.A(\round_logic.mixcolumns_block_71__N_1149[6] ), 
         .B(\round_logic.mixcolumns_block_79__N_1341[6] ), .Z(n33886)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_rep_582.init = 16'h6666;
    LUT4 i3_3_lut_4_lut_adj_384 (.A(\round_logic.mixcolumns_block_71__N_1149[6] ), 
         .B(\round_logic.mixcolumns_block_79__N_1341[6] ), .C(\round_logic.mixcolumns_block_79__N_1341[5] ), 
         .D(\enc_new_block[93] ), .Z(n8_adj_8190)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i3_3_lut_4_lut_adj_384.init = 16'h6996;
    LUT4 i1_2_lut_rep_583 (.A(\enc_new_block[53] ), .B(\enc_new_block[93] ), 
         .Z(n33887)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_rep_583.init = 16'h6666;
    LUT4 i3_3_lut_4_lut_adj_385 (.A(\enc_new_block[53] ), .B(\enc_new_block[93] ), 
         .C(\enc_new_block[92] ), .D(\round_logic.mixcolumns_block_79__N_1341[6] ), 
         .Z(n8_adj_8160)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i3_3_lut_4_lut_adj_385.init = 16'h6996;
    LUT4 i1_2_lut_rep_584 (.A(\round_logic.mixcolumns_block_79__N_1341[7] ), 
         .B(\round_logic.mixcolumns_block_71__N_1149[7] ), .Z(n33888)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_rep_584.init = 16'h6666;
    LUT4 i3_3_lut_4_lut_adj_386 (.A(\round_logic.mixcolumns_block_79__N_1341[7] ), 
         .B(\round_logic.mixcolumns_block_71__N_1149[7] ), .C(\round_logic.mixcolumns_block_79__N_1341[6] ), 
         .D(\enc_new_block[94] ), .Z(n8_adj_8193)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i3_3_lut_4_lut_adj_386.init = 16'h6996;
    LUT4 i1_2_lut_rep_585 (.A(\enc_new_block[55] ), .B(\round_logic.mixcolumns_block_79__N_1341[0] ), 
         .Z(n33889)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i1_2_lut_rep_585.init = 16'h6666;
    LUT4 i3_3_lut_4_lut_adj_387 (.A(\enc_new_block[55] ), .B(\round_logic.mixcolumns_block_79__N_1341[0] ), 
         .C(\round_logic.mixcolumns_block_71__N_1149[7] ), .D(round_key[71]), 
         .Z(n8_adj_8166)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i3_3_lut_4_lut_adj_387.init = 16'h6996;
    LUT4 i2_2_lut_3_lut_adj_388 (.A(\enc_new_block[55] ), .B(\round_logic.mixcolumns_block_79__N_1341[0] ), 
         .C(round_key[81]), .Z(n7_adj_8177)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i2_2_lut_3_lut_adj_388.init = 16'h9696;
    LUT4 i1_2_lut_rep_586 (.A(\enc_new_block[94] ), .B(\enc_new_block[54] ), 
         .Z(n33890)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_rep_586.init = 16'h6666;
    LUT4 i3_3_lut_4_lut_adj_389 (.A(\enc_new_block[94] ), .B(\enc_new_block[54] ), 
         .C(round_key[70]), .D(\round_logic.mixcolumns_block_71__N_1149[6] ), 
         .Z(n8_adj_8163)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i3_3_lut_4_lut_adj_389.init = 16'h6996;
    LUT4 i1_2_lut_rep_587 (.A(\enc_new_block[82] ), .B(\round_logic.mixcolumns_block_103__N_1101[2] ), 
         .Z(n33891)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_rep_587.init = 16'h6666;
    LUT4 i3_3_lut_4_lut_adj_390 (.A(\enc_new_block[82] ), .B(\round_logic.mixcolumns_block_103__N_1101[2] ), 
         .C(\enc_new_block[122] ), .D(\enc_new_block[42] ), .Z(n8_adj_8060)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i3_3_lut_4_lut_adj_390.init = 16'h6996;
    LUT4 i1_2_lut_rep_588 (.A(\enc_new_block[2] ), .B(\enc_new_block[122] ), 
         .Z(n33892)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_rep_588.init = 16'h6666;
    LUT4 i2_2_lut_3_lut_adj_391 (.A(\enc_new_block[2] ), .B(\enc_new_block[122] ), 
         .C(round_key[99]), .Z(n7_adj_8065)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i2_2_lut_3_lut_adj_391.init = 16'h9696;
    LUT4 i3_3_lut_4_lut_adj_392 (.A(\enc_new_block[83] ), .B(\enc_new_block[123] ), 
         .C(\enc_new_block[3] ), .D(round_key[107]), .Z(n8_adj_8075)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i3_3_lut_4_lut_adj_392.init = 16'h6996;
    LUT4 i3_3_lut_4_lut_adj_393 (.A(\enc_new_block[83] ), .B(\enc_new_block[123] ), 
         .C(n33897), .D(\enc_new_block[43] ), .Z(n8_adj_8066)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i3_3_lut_4_lut_adj_393.init = 16'h6996;
    LUT4 i1_2_lut_rep_589 (.A(\enc_new_block[124] ), .B(\enc_new_block[3] ), 
         .Z(n33893)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i1_2_lut_rep_589.init = 16'h6666;
    LUT4 i1_2_lut_rep_590 (.A(\round_logic.mixcolumns_block_103__N_1101[0] ), 
         .B(\round_logic.mixcolumns_block_111__N_1285[0] ), .Z(n33894)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i1_2_lut_rep_590.init = 16'h6666;
    LUT4 i3_2_lut_3_lut_4_lut (.A(\round_logic.mixcolumns_block_103__N_1101[0] ), 
         .B(\round_logic.mixcolumns_block_111__N_1285[0] ), .C(\enc_new_block[3] ), 
         .D(\enc_new_block[124] ), .Z(n9_adj_8078)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i3_2_lut_3_lut_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_591 (.A(\enc_new_block[0] ), .B(\enc_new_block[120] ), 
         .Z(n33895)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_rep_591.init = 16'h6666;
    LUT4 i3_3_lut_4_lut_adj_394 (.A(\enc_new_block[0] ), .B(\enc_new_block[120] ), 
         .C(\round_logic.mixcolumns_block_111__N_1285[2] ), .D(n33897), 
         .Z(n8_adj_8057)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i3_3_lut_4_lut_adj_394.init = 16'h6996;
    LUT4 i1_2_lut_rep_592 (.A(\round_logic.mixcolumns_block_111__N_1285[0] ), 
         .B(\enc_new_block[87] ), .Z(n33896)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i1_2_lut_rep_592.init = 16'h6666;
    LUT4 i3_3_lut_4_lut_adj_395 (.A(\round_logic.mixcolumns_block_111__N_1285[0] ), 
         .B(\enc_new_block[87] ), .C(round_key[113]), .D(n29077), .Z(n8_adj_8085)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i3_3_lut_4_lut_adj_395.init = 16'h6996;
    LUT4 i3_3_lut_4_lut_adj_396 (.A(\round_logic.mixcolumns_block_111__N_1285[0] ), 
         .B(\enc_new_block[87] ), .C(\enc_new_block[42] ), .D(n29105), 
         .Z(n8_adj_8091)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i3_3_lut_4_lut_adj_396.init = 16'h6996;
    LUT4 i1_2_lut_rep_593 (.A(\round_logic.mixcolumns_block_103__N_1101[0] ), 
         .B(\enc_new_block[127] ), .Z(n33897)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i1_2_lut_rep_593.init = 16'h6666;
    LUT4 i3_3_lut_4_lut_adj_397 (.A(\round_logic.mixcolumns_block_103__N_1101[0] ), 
         .B(\enc_new_block[127] ), .C(round_key[119]), .D(\enc_new_block[86] ), 
         .Z(n8_adj_8103)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i3_3_lut_4_lut_adj_397.init = 16'h6996;
    LUT4 i1_2_lut_rep_594 (.A(\enc_new_block[80] ), .B(\enc_new_block[120] ), 
         .Z(n33898)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_rep_594.init = 16'h6666;
    LUT4 i3_3_lut_4_lut_adj_398 (.A(\enc_new_block[80] ), .B(\enc_new_block[120] ), 
         .C(n33903), .D(n33899), .Z(n8_adj_8109)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i3_3_lut_4_lut_adj_398.init = 16'h6996;
    LUT4 i1_2_lut_rep_595 (.A(\round_logic.mixcolumns_block_111__N_1285[2] ), 
         .B(\round_logic.mixcolumns_block_103__N_1101[2] ), .Z(n33899)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i1_2_lut_rep_595.init = 16'h6666;
    LUT4 i2_2_lut_3_lut_adj_399 (.A(\round_logic.mixcolumns_block_111__N_1285[2] ), 
         .B(\round_logic.mixcolumns_block_103__N_1101[2] ), .C(\enc_new_block[121] ), 
         .Z(n7_adj_8084)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i2_2_lut_3_lut_adj_399.init = 16'h9696;
    LUT4 i1_2_lut_rep_596 (.A(\enc_new_block[42] ), .B(\enc_new_block[2] ), 
         .Z(n33900)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_rep_596.init = 16'h6666;
    LUT4 i2_2_lut_3_lut_4_lut_adj_400 (.A(\enc_new_block[42] ), .B(\enc_new_block[2] ), 
         .C(\round_logic.mixcolumns_block_111__N_1285[0] ), .D(\round_logic.mixcolumns_block_103__N_1101[0] ), 
         .Z(n7_adj_8074)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i2_2_lut_3_lut_4_lut_adj_400.init = 16'h6996;
    LUT4 i3_3_lut_4_lut_adj_401 (.A(\enc_new_block[42] ), .B(\enc_new_block[2] ), 
         .C(round_key[114]), .D(\round_logic.mixcolumns_block_111__N_1285[2] ), 
         .Z(n8_adj_8088)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i3_3_lut_4_lut_adj_401.init = 16'h6996;
    LUT4 i1_2_lut_rep_597 (.A(\enc_new_block[121] ), .B(\enc_new_block[81] ), 
         .Z(n33901)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_rep_597.init = 16'h6666;
    LUT4 i2_2_lut_3_lut_adj_402 (.A(\enc_new_block[121] ), .B(\enc_new_block[81] ), 
         .C(\enc_new_block[40] ), .Z(n7_adj_8071)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i2_2_lut_3_lut_adj_402.init = 16'h9696;
    LUT4 \round_key_gen.trw_2__bdd_4_lut_28839  (.A(round_key[58]), .B(n11593), 
         .C(n33866), .D(\enc_new_block[18] ), .Z(n32899)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam \round_key_gen.trw_2__bdd_4_lut_28839 .init = 16'h6996;
    LUT4 i1_2_lut_adj_403 (.A(n6364[3]), .B(n6347[1]), .Z(n1)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam i1_2_lut_adj_403.init = 16'h8888;
    LUT4 i2_2_lut_3_lut_adj_404 (.A(\enc_new_block[121] ), .B(\enc_new_block[81] ), 
         .C(round_key[97]), .Z(n7_adj_8056)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i2_2_lut_3_lut_adj_404.init = 16'h9696;
    LUT4 \round_key_gen.trw_2__bdd_3_lut_28840  (.A(\round_key_gen.trw[2] ), 
         .B(n32899), .C(n33846), .Z(n32900)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \round_key_gen.trw_2__bdd_3_lut_28840 .init = 16'hcaca;
    LUT4 round_key_56__bdd_3_lut (.A(round_key[56]), .B(n33846), .C(\block_reg[2][24] ), 
         .Z(n32910)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_56__bdd_3_lut.init = 16'h4848;
    LUT4 \round_key_gen.trw_0__bdd_4_lut_28851  (.A(round_key[56]), .B(n33868), 
         .C(n33863), .D(\enc_new_block[64] ), .Z(n32912)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam \round_key_gen.trw_0__bdd_4_lut_28851 .init = 16'h6996;
    LUT4 \round_key_gen.trw_0__bdd_3_lut_28852  (.A(\round_key_gen.trw[0] ), 
         .B(n32912), .C(n33846), .Z(n32913)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \round_key_gen.trw_0__bdd_3_lut_28852 .init = 16'hcaca;
    LUT4 i15171_3_lut (.A(n33845), .B(n33846), .C(n6364_c[1]), .Z(n20693)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i15171_3_lut.init = 16'hdcdc;
    FD1P3AX block_w3_reg__i2 (.D(n5291[1]), .SP(block_w3_we), .CK(clk_c), 
            .Q(\round_logic.mixcolumns_block_103__N_1101[2] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w3_reg__i2.GSR = "ENABLED";
    LUT4 round_key_55__bdd_3_lut (.A(round_key[55]), .B(n33846), .C(\block_reg[2][23] ), 
         .Z(n32920)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_55__bdd_3_lut.init = 16'h4848;
    PFUMX i28778 (.BLUT(n33035), .ALUT(n33034), .C0(n33847), .Z(n33036));
    FD1P3AX block_w3_reg__i3 (.D(n5291[2]), .SP(block_w3_we), .CK(clk_c), 
            .Q(\enc_new_block[2] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w3_reg__i3.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i4 (.D(n5291[3]), .SP(block_w3_we), .CK(clk_c), 
            .Q(\enc_new_block[3] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w3_reg__i4.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i5 (.D(n5291[4]), .SP(block_w3_we), .CK(clk_c), 
            .Q(\round_logic.mixcolumns_block_103__N_1101[5] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w3_reg__i5.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i6 (.D(n5291[5]), .SP(block_w3_we), .CK(clk_c), 
            .Q(\round_logic.mixcolumns_block_103__N_1101[6] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w3_reg__i6.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i7 (.D(n33239), .SP(block_w3_we), .CK(clk_c), 
            .Q(\round_logic.mixcolumns_block_103__N_1101[7] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w3_reg__i7.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i8 (.D(n5291[7]), .SP(block_w3_we), .CK(clk_c), 
            .Q(\round_logic.mixcolumns_block_103__N_1101[0] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w3_reg__i8.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i9 (.D(n33227), .SP(block_w3_we), .CK(clk_c), 
            .Q(\enc_new_block[8] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w3_reg__i9.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i10 (.D(n33221), .SP(block_w3_we), .CK(clk_c), 
            .Q(\round_logic.mixcolumns_block_79__N_1341[2] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w3_reg__i10.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i11 (.D(n5291[10]), .SP(block_w3_we), .CK(clk_c), 
            .Q(\enc_new_block[10] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w3_reg__i11.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i12 (.D(n33209), .SP(block_w3_we), .CK(clk_c), 
            .Q(\enc_new_block[11] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w3_reg__i12.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i13 (.D(n5291[12]), .SP(block_w3_we), .CK(clk_c), 
            .Q(\round_logic.mixcolumns_block_79__N_1341[5] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w3_reg__i13.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i14 (.D(n33197), .SP(block_w3_we), .CK(clk_c), 
            .Q(\round_logic.mixcolumns_block_79__N_1341[6] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w3_reg__i14.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i15 (.D(n5291[14]), .SP(block_w3_we), .CK(clk_c), 
            .Q(\round_logic.mixcolumns_block_79__N_1341[7] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w3_reg__i15.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i16 (.D(n33185), .SP(block_w3_we), .CK(clk_c), 
            .Q(\round_logic.mixcolumns_block_79__N_1341[0] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w3_reg__i16.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i17 (.D(n33176), .SP(block_w3_we), .CK(clk_c), 
            .Q(\enc_new_block[16] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w3_reg__i17.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i18 (.D(n5291[17]), .SP(block_w3_we), .CK(clk_c), 
            .Q(\enc_new_block[17] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w3_reg__i18.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i19 (.D(n33162), .SP(block_w3_we), .CK(clk_c), 
            .Q(\enc_new_block[18] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w3_reg__i19.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i20 (.D(n5291[19]), .SP(block_w3_we), .CK(clk_c), 
            .Q(\enc_new_block[19] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w3_reg__i20.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i21 (.D(n5291[20]), .SP(block_w3_we), .CK(clk_c), 
            .Q(\enc_new_block[20] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w3_reg__i21.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i22 (.D(n5291[21]), .SP(block_w3_we), .CK(clk_c), 
            .Q(\enc_new_block[21] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w3_reg__i22.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i23 (.D(n33141), .SP(block_w3_we), .CK(clk_c), 
            .Q(\enc_new_block[22] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w3_reg__i23.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i24 (.D(n33135), .SP(block_w3_we), .CK(clk_c), 
            .Q(\enc_new_block[23] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w3_reg__i24.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i25 (.D(n33126), .SP(block_w3_we), .CK(clk_c), 
            .Q(\enc_new_block[24] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w3_reg__i25.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i26 (.D(n5291[25]), .SP(block_w3_we), .CK(clk_c), 
            .Q(\enc_new_block[25] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w3_reg__i26.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i27 (.D(n33112), .SP(block_w3_we), .CK(clk_c), 
            .Q(\enc_new_block[26] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w3_reg__i27.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i28 (.D(n5291[27]), .SP(block_w3_we), .CK(clk_c), 
            .Q(\enc_new_block[27] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w3_reg__i28.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i29 (.D(n5291[28]), .SP(block_w3_we), .CK(clk_c), 
            .Q(\enc_new_block[28] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w3_reg__i29.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i30 (.D(n33093), .SP(block_w3_we), .CK(clk_c), 
            .Q(\enc_new_block[29] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w3_reg__i30.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i31 (.D(n5291[30]), .SP(block_w3_we), .CK(clk_c), 
            .Q(\enc_new_block[30] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w3_reg__i31.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i32 (.D(n33081), .SP(block_w3_we), .CK(clk_c), 
            .Q(\enc_new_block[31] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w3_reg__i32.GSR = "ENABLED";
    LUT4 new_sboxw_23__bdd_4_lut_28859 (.A(round_key[55]), .B(n29123), .C(\round_logic.mixcolumns_block_47__N_1397[0] ), 
         .D(\enc_new_block[22] ), .Z(n32922)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam new_sboxw_23__bdd_4_lut_28859.init = 16'h6996;
    LUT4 new_sboxw_23__bdd_3_lut_28860 (.A(\new_sboxw[23] ), .B(n32922), 
         .C(n33846), .Z(n32923)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam new_sboxw_23__bdd_3_lut_28860.init = 16'hcaca;
    LUT4 i27389_3_lut_4_lut (.A(\block_new_127__N_1645[69] ), .B(n33846), 
         .C(n33847), .D(n13002), .Z(n5932[69])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27389_3_lut_4_lut.init = 16'hf808;
    LUT4 round_key_54__bdd_3_lut (.A(round_key[54]), .B(n33846), .C(\block_reg[2][22] ), 
         .Z(n32934)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_54__bdd_3_lut.init = 16'h4848;
    LUT4 new_sboxw_22__bdd_4_lut_28864 (.A(round_key[54]), .B(n33870), .C(n28869), 
         .D(\enc_new_block[62] ), .Z(n32936)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam new_sboxw_22__bdd_4_lut_28864.init = 16'h6996;
    LUT4 new_sboxw_22__bdd_3_lut_28865 (.A(\new_sboxw[22] ), .B(n32936), 
         .C(n33846), .Z(n32937)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam new_sboxw_22__bdd_3_lut_28865.init = 16'hcaca;
    LUT4 round_key_53__bdd_3_lut (.A(round_key[53]), .B(n33846), .C(\block_reg[2][21] ), 
         .Z(n32940)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_53__bdd_3_lut.init = 16'h4848;
    LUT4 new_sboxw_21__bdd_4_lut (.A(round_key[53]), .B(n33855), .C(\round_logic.mixcolumns_block_47__N_1397[6] ), 
         .D(\enc_new_block[20] ), .Z(n32942)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam new_sboxw_21__bdd_4_lut.init = 16'h6996;
    LUT4 new_sboxw_21__bdd_3_lut (.A(\new_sboxw[21] ), .B(n32942), .C(n33846), 
         .Z(n32943)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam new_sboxw_21__bdd_3_lut.init = 16'hcaca;
    LUT4 round_key_52__bdd_3_lut (.A(round_key[52]), .B(n33846), .C(\block_reg[2][20] ), 
         .Z(n32949)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_52__bdd_3_lut.init = 16'h4848;
    LUT4 new_sboxw_20__bdd_4_lut (.A(round_key[52]), .B(n33854), .C(n28939), 
         .D(\enc_new_block[60] ), .Z(n32951)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam new_sboxw_20__bdd_4_lut.init = 16'h6996;
    LUT4 new_sboxw_20__bdd_3_lut (.A(\new_sboxw[20] ), .B(n32951), .C(n33846), 
         .Z(n32952)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam new_sboxw_20__bdd_3_lut.init = 16'hcaca;
    LUT4 round_key_48__bdd_3_lut (.A(round_key[48]), .B(n33846), .C(\block_reg[2][16] ), 
         .Z(n32970)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_48__bdd_3_lut.init = 16'h4848;
    LUT4 new_sboxw_16__bdd_4_lut_28894 (.A(round_key[48]), .B(n29071), .C(n33933), 
         .D(\enc_new_block[104] ), .Z(n32972)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam new_sboxw_16__bdd_4_lut_28894.init = 16'h6996;
    LUT4 new_sboxw_16__bdd_3_lut_28895 (.A(\new_sboxw[16] ), .B(n32972), 
         .C(n33846), .Z(n32973)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam new_sboxw_16__bdd_3_lut_28895.init = 16'hcaca;
    LUT4 round_key_47__bdd_3_lut (.A(round_key[47]), .B(n33846), .C(\block_reg[2][15] ), 
         .Z(n32979)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_47__bdd_3_lut.init = 16'h4848;
    LUT4 \round_key_gen.trw_23__bdd_4_lut_28902  (.A(round_key[47]), .B(n29123), 
         .C(\enc_new_block[23] ), .D(\round_logic.mixcolumns_block_39__N_1197[7] ), 
         .Z(n32981)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam \round_key_gen.trw_23__bdd_4_lut_28902 .init = 16'h6996;
    LUT4 \round_key_gen.trw_23__bdd_3_lut_28903  (.A(\round_key_gen.trw[23] ), 
         .B(n32981), .C(n33846), .Z(n32982)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \round_key_gen.trw_23__bdd_3_lut_28903 .init = 16'hcaca;
    LUT4 round_key_46__bdd_3_lut (.A(round_key[46]), .B(n33846), .C(\block_reg[2][14] ), 
         .Z(n32985)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_46__bdd_3_lut.init = 16'h4848;
    LUT4 i27387_3_lut_4_lut (.A(\block_new_127__N_1645[68] ), .B(n33846), 
         .C(n33847), .D(n13001), .Z(n5932[68])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27387_3_lut_4_lut.init = 16'hf808;
    LUT4 i27385_3_lut_4_lut (.A(\block_new_127__N_1645[67] ), .B(n33846), 
         .C(n33847), .D(n13000), .Z(n5932[67])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27385_3_lut_4_lut.init = 16'hf808;
    LUT4 \round_key_gen.trw_22__bdd_4_lut_29692  (.A(round_key[46]), .B(n11620), 
         .C(n28869), .D(\round_logic.mixcolumns_block_39__N_1197[6] ), .Z(n32987)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam \round_key_gen.trw_22__bdd_4_lut_29692 .init = 16'h6996;
    LUT4 \round_key_gen.trw_22__bdd_3_lut  (.A(\round_key_gen.trw[22] ), .B(n32987), 
         .C(n33846), .Z(n32988)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \round_key_gen.trw_22__bdd_3_lut .init = 16'hcaca;
    LUT4 round_key_45__bdd_3_lut (.A(round_key[45]), .B(n33846), .C(\block_reg[2][13] ), 
         .Z(n32994)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_45__bdd_3_lut.init = 16'h4848;
    FD1P3AX block_w0_reg__i2 (.D(n5291[97]), .SP(block_w0_we), .CK(clk_c), 
            .Q(\round_logic.mixcolumns_block_71__N_1149[2] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w0_reg__i2.GSR = "ENABLED";
    LUT4 \round_key_gen.trw_21__bdd_3_lut_28913  (.A(\round_key_gen.trw[21] ), 
         .B(n32996), .C(n33846), .Z(n32997)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \round_key_gen.trw_21__bdd_3_lut_28913 .init = 16'hcaca;
    LUT4 i27381_3_lut_4_lut (.A(\block_new_127__N_1645[65] ), .B(n33846), 
         .C(n33847), .D(n12998), .Z(n5932[65])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27381_3_lut_4_lut.init = 16'hf808;
    LUT4 round_key_42__bdd_3_lut (.A(round_key[42]), .B(n33846), .C(\block_reg[2][10] ), 
         .Z(n33011)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_42__bdd_3_lut.init = 16'h4848;
    LUT4 \round_key_gen.trw_18__bdd_4_lut_29714  (.A(round_key[42]), .B(n33864), 
         .C(n33867), .D(\enc_new_block[66] ), .Z(n33013)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam \round_key_gen.trw_18__bdd_4_lut_29714 .init = 16'h6996;
    LUT4 \round_key_gen.trw_18__bdd_3_lut  (.A(\round_key_gen.trw[18] ), .B(n33013), 
         .C(n33846), .Z(n33014)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \round_key_gen.trw_18__bdd_3_lut .init = 16'hcaca;
    LUT4 i27379_3_lut_4_lut (.A(\block_new_127__N_1645[64] ), .B(n33846), 
         .C(n33847), .D(n12997), .Z(n5932[64])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27379_3_lut_4_lut.init = 16'hf808;
    LUT4 round_key_40__bdd_3_lut (.A(round_key[40]), .B(n33846), .C(\block_reg[2][8] ), 
         .Z(n33023)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_40__bdd_3_lut.init = 16'h4848;
    LUT4 \round_key_gen.trw_16__bdd_3_lut_28936  (.A(\round_key_gen.trw[16] ), 
         .B(n33025), .C(n33846), .Z(n33026)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \round_key_gen.trw_16__bdd_3_lut_28936 .init = 16'hcaca;
    PFUMX i28767 (.BLUT(n33023), .ALUT(n33022), .C0(n33847), .Z(n33024));
    PFUMX i28758 (.BLUT(n33011), .ALUT(n33010), .C0(n33847), .Z(n33012));
    PFUMX i28744 (.BLUT(n32994), .ALUT(n32993), .C0(n33847), .Z(n32995));
    LUT4 i1_2_lut_rep_598 (.A(\enc_new_block[84] ), .B(\round_logic.mixcolumns_block_111__N_1285[5] ), 
         .Z(n33902)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_rep_598.init = 16'h6666;
    PFUMX i28738 (.BLUT(n32985), .ALUT(n32984), .C0(n33847), .Z(n32986));
    LUT4 mux_692_Mux_1_i2_4_lut (.A(\round_key_gen.trw[9] ), .B(n9_adj_8207), 
         .C(n33846), .D(n10_adj_8208), .Z(n2_adj_8209)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_1_i2_4_lut.init = 16'h3aca;
    LUT4 mux_692_Mux_2_i2_4_lut (.A(\round_key_gen.trw[10] ), .B(n7_adj_8206), 
         .C(n33846), .D(n8_adj_8210), .Z(n2_adj_8211)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_2_i2_4_lut.init = 16'h3aca;
    PFUMX i28735 (.BLUT(n32979), .ALUT(n32978), .C0(n33847), .Z(n32980));
    PFUMX i28729 (.BLUT(n32970), .ALUT(n32969), .C0(n33847), .Z(n32971));
    PFUMX i28711 (.BLUT(n32949), .ALUT(n32948), .C0(n33847), .Z(n32950));
    LUT4 i1_2_lut_3_lut (.A(\enc_new_block[84] ), .B(\round_logic.mixcolumns_block_111__N_1285[5] ), 
         .C(\enc_new_block[123] ), .Z(n28933)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_3_lut.init = 16'h9696;
    PFUMX i28705 (.BLUT(n32940), .ALUT(n32939), .C0(n33847), .Z(n32941));
    PFUMX i28702 (.BLUT(n32934), .ALUT(n32933), .C0(n33847), .Z(n32935));
    LUT4 round_key_38__bdd_3_lut (.A(round_key[38]), .B(n33846), .C(\block_reg[2][6] ), 
         .Z(n33035)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_38__bdd_3_lut.init = 16'h4848;
    LUT4 mux_692_Mux_3_i2_4_lut (.A(\round_key_gen.trw[11] ), .B(n7_adj_8205), 
         .C(n33846), .D(n8_adj_8212), .Z(n2_adj_8213)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_3_i2_4_lut.init = 16'h3aca;
    LUT4 mux_692_Mux_4_i2_4_lut (.A(\round_key_gen.trw[12] ), .B(n7_adj_8204), 
         .C(n33846), .D(n8_adj_8214), .Z(n2_adj_8215)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_4_i2_4_lut.init = 16'h3aca;
    LUT4 i2_3_lut (.A(n33845), .B(n33847), .C(n33846), .Z(n5)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(291[9:20])
    defparam i2_3_lut.init = 16'hfefe;
    LUT4 mux_692_Mux_5_i2_4_lut (.A(\round_key_gen.trw[13] ), .B(n7_adj_8203), 
         .C(n33846), .D(n8_adj_8216), .Z(n2_adj_8217)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_5_i2_4_lut.init = 16'h3aca;
    PFUMX i28692 (.BLUT(n32920), .ALUT(n32919), .C0(n33847), .Z(n32921));
    LUT4 mux_692_Mux_7_i2_4_lut (.A(\round_key_gen.trw[15] ), .B(n7_adj_8202), 
         .C(n33846), .D(n8_adj_8218), .Z(n2_adj_8219)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_7_i2_4_lut.init = 16'h3aca;
    FD1P3AX block_w0_reg__i3 (.D(n5291[98]), .SP(block_w0_we), .CK(clk_c), 
            .Q(\enc_new_block[98] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w0_reg__i3.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i4 (.D(n5291[99]), .SP(block_w0_we), .CK(clk_c), 
            .Q(\enc_new_block[99] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w0_reg__i4.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i5 (.D(n32310), .SP(block_w0_we), .CK(clk_c), 
            .Q(\round_logic.mixcolumns_block_71__N_1149[5] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w0_reg__i5.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i6 (.D(n32304), .SP(block_w0_we), .CK(clk_c), 
            .Q(\round_logic.mixcolumns_block_71__N_1149[6] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w0_reg__i6.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i7 (.D(n5291[102]), .SP(block_w0_we), .CK(clk_c), 
            .Q(\round_logic.mixcolumns_block_71__N_1149[7] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w0_reg__i7.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i8 (.D(n32295), .SP(block_w0_we), .CK(clk_c), 
            .Q(\round_logic.mixcolumns_block_71__N_1149[0] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w0_reg__i8.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i9 (.D(n32289), .SP(block_w0_we), .CK(clk_c), 
            .Q(\enc_new_block[104] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w0_reg__i9.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i10 (.D(n5291[105]), .SP(block_w0_we), .CK(clk_c), 
            .Q(\round_logic.mixcolumns_block_47__N_1397[2] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w0_reg__i10.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i11 (.D(n32280), .SP(block_w0_we), .CK(clk_c), 
            .Q(\enc_new_block[106] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w0_reg__i11.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i12 (.D(n5291[107]), .SP(block_w0_we), .CK(clk_c), 
            .Q(\enc_new_block[107] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w0_reg__i12.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i13 (.D(n5291[108]), .SP(block_w0_we), .CK(clk_c), 
            .Q(\round_logic.mixcolumns_block_47__N_1397[5] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w0_reg__i13.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i14 (.D(n32266), .SP(block_w0_we), .CK(clk_c), 
            .Q(\round_logic.mixcolumns_block_47__N_1397[6] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w0_reg__i14.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i15 (.D(n32260), .SP(block_w0_we), .CK(clk_c), 
            .Q(\round_logic.mixcolumns_block_47__N_1397[7] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w0_reg__i15.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i16 (.D(n32254), .SP(block_w0_we), .CK(clk_c), 
            .Q(\round_logic.mixcolumns_block_47__N_1397[0] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w0_reg__i16.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i17 (.D(n32248), .SP(block_w0_we), .CK(clk_c), 
            .Q(\enc_new_block[112] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w0_reg__i17.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i18 (.D(n5291[113]), .SP(block_w0_we), .CK(clk_c), 
            .Q(\enc_new_block[113] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w0_reg__i18.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i19 (.D(n5291[114]), .SP(block_w0_we), .CK(clk_c), 
            .Q(\enc_new_block[114] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w0_reg__i19.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i20 (.D(n5291[115]), .SP(block_w0_we), .CK(clk_c), 
            .Q(\enc_new_block[115] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w0_reg__i20.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i21 (.D(n5291[116]), .SP(block_w0_we), .CK(clk_c), 
            .Q(\enc_new_block[116] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w0_reg__i21.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i22 (.D(n32228), .SP(block_w0_we), .CK(clk_c), 
            .Q(\enc_new_block[117] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w0_reg__i22.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i23 (.D(n5291[118]), .SP(block_w0_we), .CK(clk_c), 
            .Q(\enc_new_block[118] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w0_reg__i23.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i24 (.D(n5291[119]), .SP(block_w0_we), .CK(clk_c), 
            .Q(\enc_new_block[119] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w0_reg__i24.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i25 (.D(n32216), .SP(block_w0_we), .CK(clk_c), 
            .Q(\enc_new_block[120] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w0_reg__i25.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i26 (.D(n5291[121]), .SP(block_w0_we), .CK(clk_c), 
            .Q(\enc_new_block[121] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w0_reg__i26.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i27 (.D(n32207), .SP(block_w0_we), .CK(clk_c), 
            .Q(\enc_new_block[122] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w0_reg__i27.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i28 (.D(n5291[123]), .SP(block_w0_we), .CK(clk_c), 
            .Q(\enc_new_block[123] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w0_reg__i28.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i29 (.D(n32198), .SP(block_w0_we), .CK(clk_c), 
            .Q(\enc_new_block[124] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w0_reg__i29.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i30 (.D(n5291[125]), .SP(block_w0_we), .CK(clk_c), 
            .Q(\enc_new_block[125] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w0_reg__i30.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i31 (.D(n32187), .SP(block_w0_we), .CK(clk_c), 
            .Q(\enc_new_block[126] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w0_reg__i31.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i32 (.D(n32181), .SP(block_w0_we), .CK(clk_c), 
            .Q(\enc_new_block[127] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w0_reg__i32.GSR = "ENABLED";
    PFUMX i28685 (.BLUT(n32910), .ALUT(n32909), .C0(n33847), .Z(n32911));
    FD1P3AX block_w1_reg__i2 (.D(n5291[65]), .SP(block_w1_we), .CK(clk_c), 
            .Q(\round_logic.mixcolumns_block_39__N_1197[2] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w1_reg__i2.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i3 (.D(n32789), .SP(block_w1_we), .CK(clk_c), 
            .Q(\enc_new_block[66] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w1_reg__i3.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i4 (.D(n5291[67]), .SP(block_w1_we), .CK(clk_c), 
            .Q(\enc_new_block[67] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w1_reg__i4.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i5 (.D(n5291[68]), .SP(block_w1_we), .CK(clk_c), 
            .Q(\round_logic.mixcolumns_block_39__N_1197[5] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w1_reg__i5.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i6 (.D(n5291[69]), .SP(block_w1_we), .CK(clk_c), 
            .Q(\round_logic.mixcolumns_block_39__N_1197[6] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w1_reg__i6.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i7 (.D(n5291[70]), .SP(block_w1_we), .CK(clk_c), 
            .Q(\round_logic.mixcolumns_block_39__N_1197[7] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w1_reg__i7.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i8 (.D(n5291[71]), .SP(block_w1_we), .CK(clk_c), 
            .Q(\round_logic.mixcolumns_block_39__N_1197[0] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w1_reg__i8.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i9 (.D(n32702), .SP(block_w1_we), .CK(clk_c), 
            .Q(\enc_new_block[72] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w1_reg__i9.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i10 (.D(n5291[73]), .SP(block_w1_we), .CK(clk_c), 
            .Q(\round_logic.mixcolumns_block_15__N_1453[2] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w1_reg__i10.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i11 (.D(n32605), .SP(block_w1_we), .CK(clk_c), 
            .Q(\enc_new_block[74] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w1_reg__i11.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i12 (.D(n5291[75]), .SP(block_w1_we), .CK(clk_c), 
            .Q(\enc_new_block[75] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w1_reg__i12.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i13 (.D(n5291[76]), .SP(block_w1_we), .CK(clk_c), 
            .Q(\round_logic.mixcolumns_block_15__N_1453[5] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w1_reg__i13.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i14 (.D(n32582), .SP(block_w1_we), .CK(clk_c), 
            .Q(\round_logic.mixcolumns_block_15__N_1453[6] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w1_reg__i14.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i15 (.D(n32576), .SP(block_w1_we), .CK(clk_c), 
            .Q(\round_logic.mixcolumns_block_15__N_1453[7] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w1_reg__i15.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i16 (.D(n32565), .SP(block_w1_we), .CK(clk_c), 
            .Q(\round_logic.mixcolumns_block_15__N_1453[0] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w1_reg__i16.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i17 (.D(n32559), .SP(block_w1_we), .CK(clk_c), 
            .Q(\enc_new_block[80] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w1_reg__i17.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i18 (.D(n5291[81]), .SP(block_w1_we), .CK(clk_c), 
            .Q(\enc_new_block[81] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w1_reg__i18.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i19 (.D(n5291[82]), .SP(block_w1_we), .CK(clk_c), 
            .Q(\enc_new_block[82] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w1_reg__i19.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i20 (.D(n5291[83]), .SP(block_w1_we), .CK(clk_c), 
            .Q(\enc_new_block[83] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w1_reg__i20.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i21 (.D(n5291[84]), .SP(block_w1_we), .CK(clk_c), 
            .Q(\enc_new_block[84] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w1_reg__i21.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i22 (.D(n5291[85]), .SP(block_w1_we), .CK(clk_c), 
            .Q(\enc_new_block[85] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w1_reg__i22.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i23 (.D(n5291[86]), .SP(block_w1_we), .CK(clk_c), 
            .Q(\enc_new_block[86] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w1_reg__i23.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i24 (.D(n5291[87]), .SP(block_w1_we), .CK(clk_c), 
            .Q(\enc_new_block[87] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w1_reg__i24.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i25 (.D(n32513), .SP(block_w1_we), .CK(clk_c), 
            .Q(\enc_new_block[88] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w1_reg__i25.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i26 (.D(n5291[89]), .SP(block_w1_we), .CK(clk_c), 
            .Q(\enc_new_block[89] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w1_reg__i26.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i27 (.D(n32367), .SP(block_w1_we), .CK(clk_c), 
            .Q(\enc_new_block[90] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w1_reg__i27.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i28 (.D(n5291[91]), .SP(block_w1_we), .CK(clk_c), 
            .Q(\enc_new_block[91] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w1_reg__i28.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i29 (.D(n5291[92]), .SP(block_w1_we), .CK(clk_c), 
            .Q(\enc_new_block[92] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w1_reg__i29.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i30 (.D(n32343), .SP(block_w1_we), .CK(clk_c), 
            .Q(\enc_new_block[93] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w1_reg__i30.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i31 (.D(n32337), .SP(block_w1_we), .CK(clk_c), 
            .Q(\enc_new_block[94] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w1_reg__i31.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i32 (.D(n32331), .SP(block_w1_we), .CK(clk_c), 
            .Q(\enc_new_block[95] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w1_reg__i32.GSR = "ENABLED";
    LUT4 mux_692_Mux_10_i2_4_lut (.A(\round_key_gen.trw[18] ), .B(n7_adj_8201), 
         .C(n33846), .D(n8_adj_8220), .Z(n2_adj_8221)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_10_i2_4_lut.init = 16'h3aca;
    LUT4 mux_692_Mux_12_i2_4_lut (.A(\round_key_gen.trw[20] ), .B(n7_adj_8222), 
         .C(n33846), .D(n8_adj_8223), .Z(n2_adj_8224)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_12_i2_4_lut.init = 16'h3aca;
    LUT4 mux_692_Mux_14_i2_4_lut (.A(\round_key_gen.trw[22] ), .B(n7_adj_8199), 
         .C(n33846), .D(n8_adj_8225), .Z(n2_adj_8226)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_14_i2_4_lut.init = 16'h3aca;
    PFUMX i28676 (.BLUT(n32897), .ALUT(n32896), .C0(n33847), .Z(n32898));
    LUT4 mux_692_Mux_17_i2_4_lut (.A(\new_sboxw[17] ), .B(n9_adj_8227), 
         .C(n33846), .D(n10_adj_8198), .Z(n2_adj_8228)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam mux_692_Mux_17_i2_4_lut.init = 16'h3aca;
    FD1P3IX round_ctr_reg_910__i3 (.D(n21[3]), .SP(round_ctr_we), .CD(n33913), 
            .CK(clk_c), .Q(enc_round_nr[3]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(387[27:47])
    defparam round_ctr_reg_910__i3.GSR = "ENABLED";
    FD1P3IX round_ctr_reg_910__i2 (.D(n21[2]), .SP(round_ctr_we), .CD(n33913), 
            .CK(clk_c), .Q(enc_round_nr[2]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(387[27:47])
    defparam round_ctr_reg_910__i2.GSR = "ENABLED";
    FD1P3IX round_ctr_reg_910__i1 (.D(n21[1]), .SP(round_ctr_we), .CD(n33913), 
            .CK(clk_c), .Q(enc_round_nr[1]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(387[27:47])
    defparam round_ctr_reg_910__i1.GSR = "ENABLED";
    FD1P3AX sword_ctr_reg_FSM_i0_i3 (.D(n28860), .SP(sword_ctr_we), .CK(clk_c), 
            .Q(n6364[3]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam sword_ctr_reg_FSM_i0_i3.GSR = "ENABLED";
    FD1P3AX sword_ctr_reg_FSM_i0_i2 (.D(n28861), .SP(sword_ctr_we), .CK(clk_c), 
            .Q(block_w2_we_N_1489));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam sword_ctr_reg_FSM_i0_i2.GSR = "ENABLED";
    FD1P3IX sword_ctr_reg_FSM_i0_i1 (.D(n6364_c[0]), .SP(sword_ctr_we), 
            .CD(n33915), .CK(clk_c), .Q(n6364_c[1]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(364[27:47])
    defparam sword_ctr_reg_FSM_i0_i1.GSR = "ENABLED";
    FD1P3IX round_ctr_reg_910__i0 (.D(n21[0]), .SP(round_ctr_we), .CD(n33913), 
            .CK(clk_c), .Q(enc_round_nr[0]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(387[27:47])
    defparam round_ctr_reg_910__i0.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_599 (.A(\enc_new_block[87] ), .B(\enc_new_block[127] ), 
         .Z(n33903)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_rep_599.init = 16'h6666;
    PFUMX i28638 (.BLUT(n32851), .ALUT(n32850), .C0(n33847), .Z(n32852));
    LUT4 i2_2_lut_3_lut_adj_405 (.A(\enc_new_block[87] ), .B(\enc_new_block[127] ), 
         .C(\enc_new_block[83] ), .Z(n7_adj_8111)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i2_2_lut_3_lut_adj_405.init = 16'h9696;
    FD1P3AX block_w2_reg__i2 (.D(n5291[33]), .SP(block_w2_we), .CK(clk_c), 
            .Q(\round_logic.mixcolumns_block_7__N_1245[2] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w2_reg__i2.GSR = "ENABLED";
    PFUMX i28589 (.BLUT(n32785), .ALUT(n32784), .C0(n33847), .Z(n32786));
    LUT4 i1_2_lut_rep_600 (.A(\enc_new_block[83] ), .B(\round_logic.mixcolumns_block_103__N_1101[5] ), 
         .Z(n33904)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i1_2_lut_rep_600.init = 16'h6666;
    FD1P3AX block_w2_reg__i3 (.D(n5291[34]), .SP(block_w2_we), .CK(clk_c), 
            .Q(\enc_new_block[34] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w2_reg__i3.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i4 (.D(n33057), .SP(block_w2_we), .CK(clk_c), 
            .Q(\enc_new_block[35] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w2_reg__i4.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i5 (.D(n5291[36]), .SP(block_w2_we), .CK(clk_c), 
            .Q(\round_logic.mixcolumns_block_7__N_1245[5] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w2_reg__i5.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i6 (.D(n5291[37]), .SP(block_w2_we), .CK(clk_c), 
            .Q(\round_logic.mixcolumns_block_7__N_1245[6] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w2_reg__i6.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i7 (.D(n33039), .SP(block_w2_we), .CK(clk_c), 
            .Q(\round_logic.mixcolumns_block_7__N_1245[7] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w2_reg__i7.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i8 (.D(n5291[39]), .SP(block_w2_we), .CK(clk_c), 
            .Q(\round_logic.mixcolumns_block_7__N_1245[0] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w2_reg__i8.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i9 (.D(n33027), .SP(block_w2_we), .CK(clk_c), 
            .Q(\enc_new_block[40] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w2_reg__i9.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i10 (.D(n5291[41]), .SP(block_w2_we), .CK(clk_c), 
            .Q(\round_logic.mixcolumns_block_111__N_1285[2] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w2_reg__i10.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i11 (.D(n33015), .SP(block_w2_we), .CK(clk_c), 
            .Q(\enc_new_block[42] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w2_reg__i11.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i12 (.D(n5291[43]), .SP(block_w2_we), .CK(clk_c), 
            .Q(\enc_new_block[43] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w2_reg__i12.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i13 (.D(n5291[44]), .SP(block_w2_we), .CK(clk_c), 
            .Q(\round_logic.mixcolumns_block_111__N_1285[5] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w2_reg__i13.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i14 (.D(n32998), .SP(block_w2_we), .CK(clk_c), 
            .Q(\round_logic.mixcolumns_block_111__N_1285[6] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w2_reg__i14.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i15 (.D(n32989), .SP(block_w2_we), .CK(clk_c), 
            .Q(\round_logic.mixcolumns_block_111__N_1285[7] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w2_reg__i15.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i16 (.D(n32983), .SP(block_w2_we), .CK(clk_c), 
            .Q(\round_logic.mixcolumns_block_111__N_1285[0] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w2_reg__i16.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i17 (.D(n32974), .SP(block_w2_we), .CK(clk_c), 
            .Q(\enc_new_block[48] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w2_reg__i17.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i18 (.D(n5291[49]), .SP(block_w2_we), .CK(clk_c), 
            .Q(\enc_new_block[49] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w2_reg__i18.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i19 (.D(n5291[50]), .SP(block_w2_we), .CK(clk_c), 
            .Q(\enc_new_block[50] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w2_reg__i19.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i20 (.D(n5291[51]), .SP(block_w2_we), .CK(clk_c), 
            .Q(\enc_new_block[51] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w2_reg__i20.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i21 (.D(n32953), .SP(block_w2_we), .CK(clk_c), 
            .Q(\enc_new_block[52] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w2_reg__i21.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i22 (.D(n32944), .SP(block_w2_we), .CK(clk_c), 
            .Q(\enc_new_block[53] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w2_reg__i22.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i23 (.D(n32938), .SP(block_w2_we), .CK(clk_c), 
            .Q(\enc_new_block[54] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w2_reg__i23.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i24 (.D(n32924), .SP(block_w2_we), .CK(clk_c), 
            .Q(\enc_new_block[55] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w2_reg__i24.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i25 (.D(n32914), .SP(block_w2_we), .CK(clk_c), 
            .Q(\enc_new_block[56] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w2_reg__i25.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i26 (.D(n5291[57]), .SP(block_w2_we), .CK(clk_c), 
            .Q(\enc_new_block[57] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w2_reg__i26.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i27 (.D(n32901), .SP(block_w2_we), .CK(clk_c), 
            .Q(\enc_new_block[58] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w2_reg__i27.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i28 (.D(n5291[59]), .SP(block_w2_we), .CK(clk_c), 
            .Q(\enc_new_block[59] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w2_reg__i28.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i29 (.D(n5291[60]), .SP(block_w2_we), .CK(clk_c), 
            .Q(\enc_new_block[60] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w2_reg__i29.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i30 (.D(n5291[61]), .SP(block_w2_we), .CK(clk_c), 
            .Q(\enc_new_block[61] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w2_reg__i30.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i31 (.D(n5291[62]), .SP(block_w2_we), .CK(clk_c), 
            .Q(\enc_new_block[62] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w2_reg__i31.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i32 (.D(n32855), .SP(block_w2_we), .CK(clk_c), 
            .Q(\enc_new_block[63] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=116, LSE_RLINE=132 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(229[9] 253[12])
    defparam block_w2_reg__i32.GSR = "ENABLED";
    LUT4 \round_key_gen.trw_16__bdd_3_lut_28937_4_lut  (.A(\enc_new_block[32] ), 
         .B(n33929), .C(n12156), .D(round_key[8]), .Z(n33225)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam \round_key_gen.trw_16__bdd_3_lut_28937_4_lut .init = 16'h6996;
    PFUMX i28523 (.BLUT(n32698), .ALUT(n32697), .C0(n33847), .Z(n32699));
    LUT4 i3_2_lut_3_lut_adj_406 (.A(\enc_new_block[83] ), .B(\round_logic.mixcolumns_block_103__N_1101[5] ), 
         .C(\enc_new_block[124] ), .Z(n9_adj_8093)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i3_2_lut_3_lut_adj_406.init = 16'h9696;
    LUT4 i1_2_lut_rep_601 (.A(\enc_new_block[124] ), .B(\round_logic.mixcolumns_block_111__N_1285[6] ), 
         .Z(n33905)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_rep_601.init = 16'h6666;
    LUT4 i3_3_lut_4_lut_adj_407 (.A(\enc_new_block[26] ), .B(n33924), .C(round_key[27]), 
         .D(\enc_new_block[114] ), .Z(n8_adj_8042)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i3_3_lut_4_lut_adj_407.init = 16'h6996;
    LUT4 i3_3_lut_4_lut_adj_408 (.A(\enc_new_block[26] ), .B(n33924), .C(\enc_new_block[34] ), 
         .D(n33922), .Z(n8_adj_8212)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i3_3_lut_4_lut_adj_408.init = 16'h6996;
    LUT4 i3_3_lut_4_lut_adj_409 (.A(\enc_new_block[64] ), .B(n33871), .C(n11593), 
         .D(\enc_new_block[104] ), .Z(n8_adj_8106)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i3_3_lut_4_lut_adj_409.init = 16'h6996;
    LUT4 \round_key_gen.trw_16__bdd_3_lut_28770_4_lut  (.A(\enc_new_block[64] ), 
         .B(n33871), .C(n33865), .D(round_key[40]), .Z(n33025)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam \round_key_gen.trw_16__bdd_3_lut_28770_4_lut .init = 16'h6996;
    LUT4 i3_3_lut_4_lut_adj_410 (.A(\enc_new_block[67] ), .B(n33871), .C(n33869), 
         .D(round_key[44]), .Z(n8_adj_8121)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i3_3_lut_4_lut_adj_410.init = 16'h6996;
    LUT4 i3_3_lut_4_lut_adj_411 (.A(\enc_new_block[67] ), .B(n33871), .C(round_key[43]), 
         .D(n33866), .Z(n8_adj_8118)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i3_3_lut_4_lut_adj_411.init = 16'h6996;
    LUT4 i3_3_lut_4_lut_adj_412 (.A(\enc_new_block[107] ), .B(n33933), .C(round_key[51]), 
         .D(\enc_new_block[18] ), .Z(n8_adj_8132)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i3_3_lut_4_lut_adj_412.init = 16'h6996;
    LUT4 \round_key_gen.trw_21__bdd_3_lut_28746_4_lut  (.A(\round_logic.mixcolumns_block_47__N_1397[5] ), 
         .B(n33934), .C(n33931), .D(round_key[45]), .Z(n32996)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam \round_key_gen.trw_21__bdd_3_lut_28746_4_lut .init = 16'h6996;
    LUT4 i3_3_lut_4_lut_adj_413 (.A(\enc_new_block[124] ), .B(\round_logic.mixcolumns_block_111__N_1285[6] ), 
         .C(round_key[125]), .D(\enc_new_block[85] ), .Z(n8_adj_8115)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i3_3_lut_4_lut_adj_413.init = 16'h6996;
    PFUMX i28446 (.BLUT(n32601), .ALUT(n32600), .C0(n33847), .Z(n32602));
    LUT4 i1_2_lut_rep_602 (.A(\enc_new_block[85] ), .B(\enc_new_block[125] ), 
         .Z(n33906)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_rep_602.init = 16'h6666;
    PFUMX i28426 (.BLUT(n32578), .ALUT(n32577), .C0(n33847), .Z(n32579));
    PFUMX i28421 (.BLUT(n32572), .ALUT(n32571), .C0(n33847), .Z(n32573));
    PFUMX i28413 (.BLUT(n32561), .ALUT(n32560), .C0(n33847), .Z(n32562));
    PFUMX i28408 (.BLUT(n32555), .ALUT(n32554), .C0(n33847), .Z(n32556));
    LUT4 i1_2_lut_rep_548_3_lut (.A(\enc_new_block[85] ), .B(\enc_new_block[125] ), 
         .C(\round_logic.mixcolumns_block_103__N_1101[5] ), .Z(n33852)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_rep_548_3_lut.init = 16'h9696;
    PFUMX i28369 (.BLUT(n32509), .ALUT(n32508), .C0(n33847), .Z(n32510));
    LUT4 i1_2_lut_rep_603 (.A(\round_logic.mixcolumns_block_111__N_1285[7] ), 
         .B(\round_logic.mixcolumns_block_103__N_1101[7] ), .Z(n33907)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_rep_603.init = 16'h6666;
    LUT4 i3_3_lut_4_lut_adj_414 (.A(\round_logic.mixcolumns_block_111__N_1285[7] ), 
         .B(\round_logic.mixcolumns_block_103__N_1101[7] ), .C(round_key[118]), 
         .D(\enc_new_block[126] ), .Z(n8_adj_8100)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i3_3_lut_4_lut_adj_414.init = 16'h6996;
    LUT4 i1_2_lut_rep_604 (.A(\enc_new_block[126] ), .B(\enc_new_block[86] ), 
         .Z(n33908)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_rep_604.init = 16'h6666;
    LUT4 \round_key_gen.trw_14__bdd_4_lut_28947  (.A(round_key[38]), .B(n11620), 
         .C(n33934), .D(\round_logic.mixcolumns_block_47__N_1397[7] ), .Z(n33037)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam \round_key_gen.trw_14__bdd_4_lut_28947 .init = 16'h6996;
    LUT4 \round_key_gen.trw_14__bdd_3_lut_28948  (.A(\round_key_gen.trw[14] ), 
         .B(n33037), .C(n33846), .Z(n33038)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \round_key_gen.trw_14__bdd_3_lut_28948 .init = 16'hcaca;
    LUT4 i27375_3_lut_4_lut (.A(\block_new_127__N_1645[62] ), .B(n33846), 
         .C(n33847), .D(n12995), .Z(n5932[62])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27375_3_lut_4_lut.init = 16'hf808;
    LUT4 i27373_3_lut_4_lut (.A(\block_new_127__N_1645[61] ), .B(n33846), 
         .C(n33847), .D(n12994), .Z(n5932[61])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27373_3_lut_4_lut.init = 16'hf808;
    LUT4 i3_3_lut_4_lut_adj_415 (.A(\enc_new_block[126] ), .B(\enc_new_block[86] ), 
         .C(\round_logic.mixcolumns_block_103__N_1101[6] ), .D(\round_logic.mixcolumns_block_111__N_1285[7] ), 
         .Z(n8_adj_8069)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i3_3_lut_4_lut_adj_415.init = 16'h6996;
    LUT4 i1_2_lut_rep_558 (.A(\round_logic.mixcolumns_block_39__N_1197[0] ), 
         .B(\enc_new_block[63] ), .Z(n33862)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i1_2_lut_rep_558.init = 16'h6666;
    LUT4 i3_3_lut_4_lut_adj_416 (.A(\round_logic.mixcolumns_block_39__N_1197[0] ), 
         .B(\enc_new_block[63] ), .C(n33869), .D(n33932), .Z(n8_adj_8063)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i3_3_lut_4_lut_adj_416.init = 16'h6996;
    LUT4 i3_3_lut_4_lut_adj_417 (.A(\round_logic.mixcolumns_block_39__N_1197[0] ), 
         .B(\enc_new_block[63] ), .C(n11593), .D(n29071), .Z(n8_adj_8051)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i3_3_lut_4_lut_adj_417.init = 16'h6996;
    LUT4 i1_2_lut_3_lut_adj_418 (.A(\round_logic.mixcolumns_block_39__N_1197[0] ), 
         .B(\enc_new_block[63] ), .C(\round_logic.mixcolumns_block_47__N_1397[7] ), 
         .Z(n29123)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i1_2_lut_3_lut_adj_418.init = 16'h9696;
    LUT4 i1_2_lut_rep_559 (.A(\enc_new_block[104] ), .B(\enc_new_block[16] ), 
         .Z(n33863)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i1_2_lut_rep_559.init = 16'h6666;
    LUT4 i3_3_lut_4_lut_adj_419 (.A(\enc_new_block[104] ), .B(\enc_new_block[16] ), 
         .C(\enc_new_block[57] ), .D(n33864), .Z(n8_adj_8126)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i3_3_lut_4_lut_adj_419.init = 16'h6996;
    LUT4 i1_2_lut_rep_560 (.A(\round_logic.mixcolumns_block_47__N_1397[2] ), 
         .B(\round_logic.mixcolumns_block_39__N_1197[2] ), .Z(n33864)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_rep_560.init = 16'h6666;
    LUT4 i2_2_lut_3_lut_adj_420 (.A(\round_logic.mixcolumns_block_47__N_1397[2] ), 
         .B(\round_logic.mixcolumns_block_39__N_1197[2] ), .C(round_key[57]), 
         .Z(n7_adj_8134)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i2_2_lut_3_lut_adj_420.init = 16'h9696;
    LUT4 i1_2_lut_rep_561 (.A(\enc_new_block[16] ), .B(\enc_new_block[56] ), 
         .Z(n33865)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_rep_561.init = 16'h6666;
    LUT4 i3_3_lut_4_lut_adj_421 (.A(\enc_new_block[16] ), .B(\enc_new_block[56] ), 
         .C(n33868), .D(\enc_new_block[17] ), .Z(n8_adj_8135)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i3_3_lut_4_lut_adj_421.init = 16'h6996;
    LUT4 i1_2_lut_rep_562 (.A(\enc_new_block[66] ), .B(\enc_new_block[106] ), 
         .Z(n33866)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_rep_562.init = 16'h6666;
    LUT4 i3_3_lut_4_lut_adj_422 (.A(\enc_new_block[66] ), .B(\enc_new_block[106] ), 
         .C(\round_logic.mixcolumns_block_47__N_1397[2] ), .D(round_key[50]), 
         .Z(n8_adj_8129)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i3_3_lut_4_lut_adj_422.init = 16'h6996;
    LUT4 i2_2_lut_adj_423 (.A(\enc_new_block[85] ), .B(\round_logic.mixcolumns_block_111__N_1285[6] ), 
         .Z(n7_adj_8099)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i2_2_lut_adj_423.init = 16'h6666;
    LUT4 i20145_3_lut_4_lut (.A(enc_round_nr[1]), .B(enc_round_nr[0]), .C(enc_round_nr[2]), 
         .D(enc_round_nr[3]), .Z(n21[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(387[27:47])
    defparam i20145_3_lut_4_lut.init = 16'h7f80;
    LUT4 i20138_2_lut_3_lut (.A(enc_round_nr[1]), .B(enc_round_nr[0]), .C(enc_round_nr[2]), 
         .Z(n21[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(387[27:47])
    defparam i20138_2_lut_3_lut.init = 16'h7878;
    LUT4 i9395_4_lut_3_lut_rep_610 (.A(enc_round_nr[2]), .B(enc_round_nr[1]), 
         .C(\key_mem_ctrl.num_rounds[2] ), .Z(n33914)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;
    defparam i9395_4_lut_3_lut_rep_610.init = 16'h8e8e;
    LUT4 i1_2_lut_rep_544_4_lut (.A(enc_round_nr[2]), .B(enc_round_nr[1]), 
         .C(\key_mem_ctrl.num_rounds[2] ), .D(enc_round_nr[3]), .Z(n33848)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A !((C+!(D))+!B)) */ ;
    defparam i1_2_lut_rep_544_4_lut.init = 16'h8e00;
    LUT4 i1_2_lut_4_lut (.A(enc_round_nr[2]), .B(enc_round_nr[1]), .C(\key_mem_ctrl.num_rounds[2] ), 
         .D(n6347[0]), .Z(n4)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A !((C+!(D))+!B)) */ ;
    defparam i1_2_lut_4_lut.init = 16'h8e00;
    LUT4 i1_2_lut_rep_611 (.A(n6347[0]), .B(n6347[2]), .Z(n33915)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(422[7] 479[14])
    defparam i1_2_lut_rep_611.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n6347[0]), .B(n6347[2]), .C(block_w2_we_N_1489), 
         .D(n6347[1]), .Z(n28860)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(422[7] 479[14])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_424 (.A(n6347[0]), .B(n6347[2]), .C(n6364_c[1]), 
         .D(n6347[1]), .Z(n28861)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(422[7] 479[14])
    defparam i1_2_lut_3_lut_4_lut_adj_424.init = 16'h1000;
    LUT4 i2_3_lut_4_lut (.A(n6347[0]), .B(n6347[2]), .C(n33913), .D(n1), 
         .Z(enc_ctrl_we)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(422[7] 479[14])
    defparam i2_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_adj_425 (.A(n6347[0]), .B(n6347[2]), .C(n6347[1]), 
         .Z(sword_ctr_we)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(422[7] 479[14])
    defparam i1_2_lut_3_lut_adj_425.init = 16'hfefe;
    LUT4 i2_3_lut_4_lut_adj_426 (.A(n6347[0]), .B(n6347[2]), .C(n6364[3]), 
         .D(n6347[1]), .Z(n25323)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(422[7] 479[14])
    defparam i2_3_lut_4_lut_adj_426.init = 16'hfeff;
    LUT4 i1_2_lut_rep_613 (.A(\round_logic.mixcolumns_block_7__N_1245[2] ), 
         .B(\enc_new_block[72] ), .Z(n33917)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i1_2_lut_rep_613.init = 16'h6666;
    LUT4 i1_2_lut_adj_427 (.A(\round_logic.mixcolumns_block_111__N_1285[6] ), 
         .B(\round_logic.mixcolumns_block_103__N_1101[6] ), .Z(n29303)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_adj_427.init = 16'h6666;
    LUT4 i1_2_lut_rep_614 (.A(\enc_new_block[26] ), .B(\round_logic.mixcolumns_block_15__N_1453[2] ), 
         .Z(n33918)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_rep_614.init = 16'h6666;
    LUT4 i4_4_lut_adj_428 (.A(\round_logic.mixcolumns_block_111__N_1285[5] ), 
         .B(round_key[116]), .C(n33896), .D(\enc_new_block[43] ), .Z(n10_adj_8094)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i4_4_lut_adj_428.init = 16'h6996;
    LUT4 i3_3_lut_4_lut_adj_429 (.A(\enc_new_block[26] ), .B(\round_logic.mixcolumns_block_15__N_1453[2] ), 
         .C(\enc_new_block[34] ), .D(round_key[10]), .Z(n8_adj_8220)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i3_3_lut_4_lut_adj_429.init = 16'h6996;
    LUT4 i2_2_lut_3_lut_adj_430 (.A(\enc_new_block[114] ), .B(\enc_new_block[74] ), 
         .C(round_key[19]), .Z(n7)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i2_2_lut_3_lut_adj_430.init = 16'h9696;
    LUT4 i3_3_lut_4_lut_adj_431 (.A(\enc_new_block[114] ), .B(\enc_new_block[74] ), 
         .C(\enc_new_block[26] ), .D(\round_logic.mixcolumns_block_7__N_1245[2] ), 
         .Z(n8_adj_8210)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i3_3_lut_4_lut_adj_431.init = 16'h6996;
    LUT4 i3_3_lut_4_lut_adj_432 (.A(\enc_new_block[35] ), .B(\enc_new_block[75] ), 
         .C(\enc_new_block[27] ), .D(n33920), .Z(n8)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i3_3_lut_4_lut_adj_432.init = 16'h6996;
    LUT4 i3_3_lut_4_lut_adj_433 (.A(\enc_new_block[35] ), .B(\enc_new_block[75] ), 
         .C(n11634), .D(\round_logic.mixcolumns_block_7__N_1245[5] ), .Z(n8_adj_8223)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i3_3_lut_4_lut_adj_433.init = 16'h6996;
    LUT4 i1_2_lut_rep_615 (.A(\round_logic.mixcolumns_block_7__N_1245[5] ), 
         .B(\round_logic.mixcolumns_block_15__N_1453[5] ), .Z(n33919)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_rep_615.init = 16'h6666;
    LUT4 i2_2_lut_3_lut_adj_434 (.A(\round_logic.mixcolumns_block_7__N_1245[5] ), 
         .B(\round_logic.mixcolumns_block_15__N_1453[5] ), .C(round_key[20]), 
         .Z(n7_adj_8025)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i2_2_lut_3_lut_adj_434.init = 16'h9696;
    LUT4 i1_2_lut_rep_616 (.A(\round_logic.mixcolumns_block_15__N_1453[0] ), 
         .B(\enc_new_block[119] ), .Z(n33920)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i1_2_lut_rep_616.init = 16'h6666;
    LUT4 i3_3_lut_4_lut_adj_435 (.A(\round_logic.mixcolumns_block_15__N_1453[0] ), 
         .B(\enc_new_block[119] ), .C(\enc_new_block[28] ), .D(n33924), 
         .Z(n8_adj_8026)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i3_3_lut_4_lut_adj_435.init = 16'h6996;
    LUT4 i2_2_lut_adj_436 (.A(\enc_new_block[123] ), .B(round_key[115]), 
         .Z(n7_adj_8090)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i2_2_lut_adj_436.init = 16'h6666;
    LUT4 i3_3_lut_4_lut_adj_437 (.A(\round_logic.mixcolumns_block_15__N_1453[0] ), 
         .B(\enc_new_block[119] ), .C(\round_logic.mixcolumns_block_7__N_1245[7] ), 
         .D(round_key[7]), .Z(n8_adj_8218)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i3_3_lut_4_lut_adj_437.init = 16'h6996;
    LUT4 i1_2_lut_rep_617 (.A(\round_logic.mixcolumns_block_7__N_1245[6] ), 
         .B(\enc_new_block[29] ), .Z(n33921)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_rep_617.init = 16'h6666;
    PFUMX i28282 (.BLUT(n32363), .ALUT(n32362), .C0(n33847), .Z(n32364));
    LUT4 i3_3_lut_4_lut_adj_438 (.A(\round_logic.mixcolumns_block_7__N_1245[6] ), 
         .B(\enc_new_block[29] ), .C(\round_logic.mixcolumns_block_15__N_1453[6] ), 
         .D(round_key[21]), .Z(n8_adj_8029)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i3_3_lut_4_lut_adj_438.init = 16'h6996;
    LUT4 i1_2_lut_rep_618 (.A(\round_logic.mixcolumns_block_7__N_1245[0] ), 
         .B(\enc_new_block[31] ), .Z(n33922)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_rep_618.init = 16'h6666;
    LUT4 i2_2_lut_adj_439 (.A(\enc_new_block[81] ), .B(\enc_new_block[122] ), 
         .Z(n7_adj_8087)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i2_2_lut_adj_439.init = 16'h6666;
    LUT4 i1_2_lut_3_lut_adj_440 (.A(\round_logic.mixcolumns_block_7__N_1245[0] ), 
         .B(\enc_new_block[31] ), .C(\round_logic.mixcolumns_block_15__N_1453[7] ), 
         .Z(n28930)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_3_lut_adj_440.init = 16'h9696;
    LUT4 i3_3_lut_4_lut_adj_441 (.A(\round_logic.mixcolumns_block_7__N_1245[0] ), 
         .B(\enc_new_block[31] ), .C(n11634), .D(n33925), .Z(n8_adj_8214)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i3_3_lut_4_lut_adj_441.init = 16'h6996;
    LUT4 i1_2_lut_rep_619 (.A(\enc_new_block[119] ), .B(\enc_new_block[112] ), 
         .Z(n33923)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i1_2_lut_rep_619.init = 16'h6666;
    LUT4 i3_2_lut_3_lut_4_lut_adj_442 (.A(\enc_new_block[119] ), .B(\enc_new_block[112] ), 
         .C(\enc_new_block[72] ), .D(\round_logic.mixcolumns_block_7__N_1245[2] ), 
         .Z(n9_adj_8227)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i3_2_lut_3_lut_4_lut_adj_442.init = 16'h6996;
    LUT4 i27275_3_lut_4_lut (.A(\block_new_127__N_1645[12] ), .B(n33846), 
         .C(n33847), .D(n12945), .Z(n5932[12])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27275_3_lut_4_lut.init = 16'hf808;
    LUT4 i1_2_lut_rep_620 (.A(\enc_new_block[75] ), .B(\enc_new_block[115] ), 
         .Z(n33924)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i1_2_lut_rep_620.init = 16'h6666;
    LUT4 i1_2_lut_adj_443 (.A(\round_logic.mixcolumns_block_103__N_1101[7] ), 
         .B(\enc_new_block[126] ), .Z(n29037)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_adj_443.init = 16'h6666;
    LUT4 i1_2_lut_rep_621 (.A(\enc_new_block[27] ), .B(\round_logic.mixcolumns_block_15__N_1453[5] ), 
         .Z(n33925)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i1_2_lut_rep_621.init = 16'h6666;
    LUT4 i27371_3_lut_4_lut (.A(\block_new_127__N_1645[60] ), .B(n33846), 
         .C(n33847), .D(n12993), .Z(n5932[60])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27371_3_lut_4_lut.init = 16'hf808;
    LUT4 i1_2_lut_rep_622 (.A(\enc_new_block[119] ), .B(\enc_new_block[31] ), 
         .Z(n33926)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i1_2_lut_rep_622.init = 16'h6666;
    LUT4 i4_4_lut_adj_444 (.A(round_key[108]), .B(\round_logic.mixcolumns_block_103__N_1101[5] ), 
         .C(\enc_new_block[84] ), .D(\enc_new_block[43] ), .Z(n10_adj_8079)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i4_4_lut_adj_444.init = 16'h6996;
    LUT4 i2_2_lut_3_lut_adj_445 (.A(\enc_new_block[119] ), .B(\enc_new_block[31] ), 
         .C(\enc_new_block[35] ), .Z(n7_adj_8041)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i2_2_lut_3_lut_adj_445.init = 16'h9696;
    LUT4 i27271_3_lut_4_lut (.A(\block_new_127__N_1645[10] ), .B(n33846), 
         .C(n33847), .D(n12943), .Z(n5932[10])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27271_3_lut_4_lut.init = 16'hf808;
    LUT4 i3_2_lut_3_lut_4_lut_adj_446 (.A(\enc_new_block[119] ), .B(\enc_new_block[31] ), 
         .C(\round_logic.mixcolumns_block_15__N_1453[5] ), .D(\enc_new_block[27] ), 
         .Z(n9_adj_8044)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i3_2_lut_3_lut_4_lut_adj_446.init = 16'h6996;
    LUT4 i27265_3_lut_4_lut (.A(\block_new_127__N_1645[7] ), .B(n33846), 
         .C(n33847), .D(n12940), .Z(n5932[7])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27265_3_lut_4_lut.init = 16'hf808;
    LUT4 i1_2_lut_rep_623 (.A(\enc_new_block[117] ), .B(\round_logic.mixcolumns_block_15__N_1453[6] ), 
         .Z(n33927)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_rep_623.init = 16'h6666;
    LUT4 i27369_3_lut_4_lut (.A(\block_new_127__N_1645[59] ), .B(n33846), 
         .C(n33847), .D(n12992), .Z(n5932[59])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27369_3_lut_4_lut.init = 16'hf808;
    LUT4 i3_3_lut_4_lut_adj_447 (.A(\enc_new_block[117] ), .B(\round_logic.mixcolumns_block_15__N_1453[6] ), 
         .C(\enc_new_block[29] ), .D(\round_logic.mixcolumns_block_7__N_1245[5] ), 
         .Z(n8_adj_8216)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i3_3_lut_4_lut_adj_447.init = 16'h6996;
    LUT4 i27261_3_lut_4_lut (.A(\block_new_127__N_1645[5] ), .B(n33846), 
         .C(n33847), .D(n12938), .Z(n5932[5])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27261_3_lut_4_lut.init = 16'hf808;
    LUT4 i27259_3_lut_4_lut (.A(\block_new_127__N_1645[4] ), .B(n33846), 
         .C(n33847), .D(n12937), .Z(n5932[4])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27259_3_lut_4_lut.init = 16'hf808;
    LUT4 i1_2_lut_rep_624 (.A(\round_logic.mixcolumns_block_7__N_1245[7] ), 
         .B(\round_logic.mixcolumns_block_15__N_1453[7] ), .Z(n33928)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_rep_624.init = 16'h6666;
    LUT4 i3_3_lut_4_lut_adj_448 (.A(\round_logic.mixcolumns_block_7__N_1245[7] ), 
         .B(\round_logic.mixcolumns_block_15__N_1453[7] ), .C(\enc_new_block[118] ), 
         .D(\enc_new_block[29] ), .Z(n8_adj_8048)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i3_3_lut_4_lut_adj_448.init = 16'h6996;
    LUT4 i1_2_lut_rep_625 (.A(\round_logic.mixcolumns_block_7__N_1245[0] ), 
         .B(\round_logic.mixcolumns_block_15__N_1453[0] ), .Z(n33929)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i1_2_lut_rep_625.init = 16'h6666;
    LUT4 i27365_3_lut_4_lut (.A(\block_new_127__N_1645[57] ), .B(n33846), 
         .C(n33847), .D(n12990), .Z(n5932[57])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27365_3_lut_4_lut.init = 16'hf808;
    LUT4 i1_2_lut_rep_549_3_lut (.A(\round_logic.mixcolumns_block_7__N_1245[0] ), 
         .B(\round_logic.mixcolumns_block_15__N_1453[0] ), .C(\enc_new_block[32] ), 
         .Z(n33853)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i1_2_lut_rep_549_3_lut.init = 16'h9696;
    LUT4 i2_2_lut_adj_449 (.A(\enc_new_block[125] ), .B(round_key[102]), 
         .Z(n7_adj_8068)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i2_2_lut_adj_449.init = 16'h6666;
    LUT4 i2_2_lut_3_lut_adj_450 (.A(\round_logic.mixcolumns_block_7__N_1245[0] ), 
         .B(\round_logic.mixcolumns_block_15__N_1453[0] ), .C(round_key[12]), 
         .Z(n7_adj_8222)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i2_2_lut_3_lut_adj_450.init = 16'h9696;
    PFUMX mux_691_i126 (.BLUT(n2_adj_8116), .ALUT(n5932[125]), .C0(n33843), 
          .Z(n5291[125]));
    LUT4 \round_key_gen.trw_19__bdd_3_lut_28923_4_lut  (.A(\round_logic.mixcolumns_block_7__N_1245[0] ), 
         .B(\round_logic.mixcolumns_block_15__N_1453[0] ), .C(n10_adj_8200), 
         .D(round_key[11]), .Z(n33207)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam \round_key_gen.trw_19__bdd_3_lut_28923_4_lut .init = 16'h6996;
    LUT4 i1_2_lut_rep_626 (.A(\enc_new_block[30] ), .B(\enc_new_block[118] ), 
         .Z(n33930)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_rep_626.init = 16'h6666;
    LUT4 i3_3_lut_4_lut_adj_451 (.A(\enc_new_block[30] ), .B(\enc_new_block[118] ), 
         .C(round_key[14]), .D(\round_logic.mixcolumns_block_7__N_1245[6] ), 
         .Z(n8_adj_8225)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i3_3_lut_4_lut_adj_451.init = 16'h6996;
    PFUMX mux_691_i124 (.BLUT(n2_adj_8113), .ALUT(n5932[123]), .C0(n33843), 
          .Z(n5291[123]));
    LUT4 i1_2_lut_rep_627 (.A(\round_logic.mixcolumns_block_39__N_1197[5] ), 
         .B(\enc_new_block[21] ), .Z(n33931)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_rep_627.init = 16'h6666;
    LUT4 i3_3_lut_4_lut_adj_452 (.A(\round_logic.mixcolumns_block_39__N_1197[5] ), 
         .B(\enc_new_block[21] ), .C(\enc_new_block[61] ), .D(\round_logic.mixcolumns_block_47__N_1397[6] ), 
         .Z(n8_adj_8082)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i3_3_lut_4_lut_adj_452.init = 16'h6996;
    LUT4 i2_2_lut_adj_453 (.A(\enc_new_block[121] ), .B(round_key[98]), 
         .Z(n7_adj_8059)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i2_2_lut_adj_453.init = 16'h6666;
    LUT4 i1_2_lut_rep_628 (.A(\enc_new_block[67] ), .B(\enc_new_block[59] ), 
         .Z(n33932)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i1_2_lut_rep_628.init = 16'h6666;
    LUT4 i2_2_lut_3_lut_adj_454 (.A(\enc_new_block[67] ), .B(\enc_new_block[59] ), 
         .C(\enc_new_block[106] ), .Z(n7_adj_8131)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i2_2_lut_3_lut_adj_454.init = 16'h9696;
    LUT4 round_key_32__bdd_3_lut (.A(round_key[32]), .B(n33846), .C(\block_reg[2][0] ), 
         .Z(n33068)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_32__bdd_3_lut.init = 16'h4848;
    PFUMX mux_691_i122 (.BLUT(n2_adj_8110), .ALUT(n5932[121]), .C0(n33843), 
          .Z(n5291[121]));
    LUT4 i1_2_lut_rep_629 (.A(\enc_new_block[23] ), .B(\round_logic.mixcolumns_block_47__N_1397[0] ), 
         .Z(n33933)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i1_2_lut_rep_629.init = 16'h6666;
    LUT4 i1_2_lut_rep_550_3_lut (.A(\enc_new_block[23] ), .B(\round_logic.mixcolumns_block_47__N_1397[0] ), 
         .C(\enc_new_block[107] ), .Z(n33854)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i1_2_lut_rep_550_3_lut.init = 16'h9696;
    LUT4 i2_2_lut_3_lut_adj_455 (.A(\enc_new_block[23] ), .B(\round_logic.mixcolumns_block_47__N_1397[0] ), 
         .C(round_key[49]), .Z(n7_adj_8125)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i2_2_lut_3_lut_adj_455.init = 16'h9696;
    PFUMX mux_691_i120 (.BLUT(n2_adj_8104), .ALUT(n5932[119]), .C0(n33843), 
          .Z(n5291[119]));
    LUT4 i3_3_lut_4_lut_adj_456 (.A(\enc_new_block[23] ), .B(\round_logic.mixcolumns_block_47__N_1397[0] ), 
         .C(\round_logic.mixcolumns_block_39__N_1197[7] ), .D(round_key[39]), 
         .Z(n8_adj_8097)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i3_3_lut_4_lut_adj_456.init = 16'h6996;
    PFUMX mux_691_i119 (.BLUT(n2_adj_8101), .ALUT(n5932[118]), .C0(n33843), 
          .Z(n5291[118]));
    LUT4 i1_2_lut_rep_630 (.A(\round_logic.mixcolumns_block_39__N_1197[6] ), 
         .B(\enc_new_block[61] ), .Z(n33934)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_rep_630.init = 16'h6666;
    LUT4 i1_2_lut_rep_551_3_lut (.A(\round_logic.mixcolumns_block_39__N_1197[6] ), 
         .B(\enc_new_block[61] ), .C(\round_logic.mixcolumns_block_47__N_1397[5] ), 
         .Z(n33855)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_rep_551_3_lut.init = 16'h9696;
    PFUMX mux_691_i117 (.BLUT(n2_adj_8095), .ALUT(n5932[116]), .C0(n33843), 
          .Z(n5291[116]));
    LUT4 i2_2_lut_adj_457 (.A(\enc_new_block[88] ), .B(round_key[89]), .Z(n7_adj_8032)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i2_2_lut_adj_457.init = 16'h6666;
    LUT4 i2_3_lut_adj_458 (.A(\enc_new_block[48] ), .B(\round_logic.mixcolumns_block_71__N_1149[2] ), 
         .C(\round_logic.mixcolumns_block_79__N_1341[2] ), .Z(n29083)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i2_3_lut_adj_458.init = 16'h9696;
    PFUMX mux_691_i116 (.BLUT(n2_adj_8092), .ALUT(n5932[115]), .C0(n33843), 
          .Z(n5291[115]));
    PFUMX mux_691_i115 (.BLUT(n2_adj_8089), .ALUT(n5932[114]), .C0(n33843), 
          .Z(n5291[114]));
    PFUMX mux_691_i114 (.BLUT(n2_adj_8086), .ALUT(n5932[113]), .C0(n33843), 
          .Z(n5291[113]));
    LUT4 i1_2_lut_adj_459 (.A(\enc_new_block[8] ), .B(\enc_new_block[96] ), 
         .Z(n29058)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_adj_459.init = 16'h6666;
    LUT4 i2_2_lut_adj_460 (.A(\round_logic.mixcolumns_block_79__N_1341[0] ), 
         .B(round_key[87]), .Z(n7_adj_8195)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i2_2_lut_adj_460.init = 16'h6666;
    LUT4 i2_2_lut_adj_461 (.A(round_key[86]), .B(\enc_new_block[53] ), .Z(n7_adj_8192)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i2_2_lut_adj_461.init = 16'h6666;
    LUT4 \round_key_gen.trw_8__bdd_4_lut_28977  (.A(round_key[32]), .B(n33862), 
         .C(n33865), .D(\enc_new_block[104] ), .Z(n33070)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam \round_key_gen.trw_8__bdd_4_lut_28977 .init = 16'h6996;
    LUT4 i2_2_lut_adj_462 (.A(round_key[85]), .B(\enc_new_block[52] ), .Z(n7_adj_8189)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i2_2_lut_adj_462.init = 16'h6666;
    LUT4 i2_2_lut_adj_463 (.A(\enc_new_block[92] ), .B(round_key[84]), .Z(n7_adj_8186)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i2_2_lut_adj_463.init = 16'h6666;
    LUT4 i2_2_lut_adj_464 (.A(round_key[82]), .B(\enc_new_block[10] ), .Z(n7_adj_8180)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i2_2_lut_adj_464.init = 16'h6666;
    LUT4 \round_key_gen.trw_8__bdd_3_lut_28978  (.A(\round_key_gen.trw[8] ), 
         .B(n33070), .C(n33846), .Z(n33071)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \round_key_gen.trw_8__bdd_3_lut_28978 .init = 16'hcaca;
    LUT4 i3_3_lut (.A(n29083), .B(\enc_new_block[8] ), .C(\enc_new_block[89] ), 
         .Z(n8_adj_8178)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i3_3_lut.init = 16'h9696;
    PFUMX mux_691_i109 (.BLUT(n2_adj_8080), .ALUT(n5932[108]), .C0(n33843), 
          .Z(n5291[108]));
    PFUMX mux_691_i108 (.BLUT(n2_adj_8076), .ALUT(n5932[107]), .C0(n33843), 
          .Z(n5291[107]));
    LUT4 round_key_31__bdd_3_lut (.A(round_key[31]), .B(n33846), .C(\block_reg[3][31] ), 
         .Z(n33077)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_31__bdd_3_lut.init = 16'h4848;
    PFUMX mux_691_i106 (.BLUT(n2_adj_8073), .ALUT(n5932[105]), .C0(n33843), 
          .Z(n5291[105]));
    PFUMX mux_691_i103 (.BLUT(n2_adj_8070), .ALUT(n5932[102]), .C0(n33843), 
          .Z(n5291[102]));
    LUT4 i2_2_lut_adj_465 (.A(\enc_new_block[95] ), .B(\enc_new_block[94] ), 
         .Z(n7_adj_8165)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i2_2_lut_adj_465.init = 16'h6666;
    LUT4 i2_2_lut_adj_466 (.A(\round_logic.mixcolumns_block_79__N_1341[7] ), 
         .B(\enc_new_block[93] ), .Z(n7_adj_8162)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i2_2_lut_adj_466.init = 16'h6666;
    LUT4 i2_2_lut_adj_467 (.A(round_key[69]), .B(\round_logic.mixcolumns_block_71__N_1149[5] ), 
         .Z(n7_adj_8159)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i2_2_lut_adj_467.init = 16'h6666;
    LUT4 i4_4_lut_adj_468 (.A(\enc_new_block[11] ), .B(\enc_new_block[90] ), 
         .C(n33877), .D(round_key[67]), .Z(n10_adj_8154)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i4_4_lut_adj_468.init = 16'h6996;
    PFUMX mux_691_i100 (.BLUT(n2_adj_8067), .ALUT(n5932[99]), .C0(n33843), 
          .Z(n5291[99]));
    PFUMX mux_691_i99 (.BLUT(n2_adj_8061), .ALUT(n5932[98]), .C0(n33843), 
          .Z(n5291[98]));
    PFUMX mux_691_i98 (.BLUT(n2_adj_8058), .ALUT(n5932[97]), .C0(n33843), 
          .Z(n5291[97]));
    PFUMX i28265 (.BLUT(n32339), .ALUT(n32338), .C0(n33847), .Z(n32340));
    LUT4 i2_2_lut_adj_469 (.A(\enc_new_block[8] ), .B(\enc_new_block[88] ), 
         .Z(n7_adj_8147)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i2_2_lut_adj_469.init = 16'h6666;
    PFUMX i28260 (.BLUT(n32333), .ALUT(n32332), .C0(n33847), .Z(n32334));
    LUT4 \round_key_gen.trw_7__bdd_4_lut_29779  (.A(round_key[31]), .B(n33929), 
         .C(n33930), .D(\enc_new_block[119] ), .Z(n33079)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam \round_key_gen.trw_7__bdd_4_lut_29779 .init = 16'h6996;
    PFUMX mux_691_i93 (.BLUT(n2_adj_8040), .ALUT(n5932[92]), .C0(n33843), 
          .Z(n5291[92]));
    LUT4 i1_2_lut_adj_470 (.A(\enc_new_block[62] ), .B(\enc_new_block[22] ), 
         .Z(n11620)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_adj_470.init = 16'h6666;
    LUT4 \round_key_gen.trw_7__bdd_3_lut  (.A(\round_key_gen.trw[7] ), .B(n33079), 
         .C(n33846), .Z(n33080)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \round_key_gen.trw_7__bdd_3_lut .init = 16'hcaca;
    LUT4 i2_2_lut_adj_471 (.A(round_key[62]), .B(\round_logic.mixcolumns_block_39__N_1197[7] ), 
         .Z(n7_adj_8144)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i2_2_lut_adj_471.init = 16'h6666;
    LUT4 round_key_29__bdd_3_lut (.A(round_key[29]), .B(n33846), .C(\block_reg[3][29] ), 
         .Z(n33089)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_29__bdd_3_lut.init = 16'h4848;
    PFUMX i28255 (.BLUT(n32327), .ALUT(n32326), .C0(n33847), .Z(n32328));
    PFUMX mux_691_i92 (.BLUT(n2_adj_8037), .ALUT(n5932[91]), .C0(n33843), 
          .Z(n5291[91]));
    LUT4 i2_2_lut_adj_472 (.A(\enc_new_block[21] ), .B(\round_logic.mixcolumns_block_47__N_1397[6] ), 
         .Z(n7_adj_8141)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i2_2_lut_adj_472.init = 16'h6666;
    LUT4 i2_2_lut_adj_473 (.A(round_key[60]), .B(\enc_new_block[20] ), .Z(n7_adj_8139)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i2_2_lut_adj_473.init = 16'h6666;
    LUT4 i2_3_lut_adj_474 (.A(\round_logic.mixcolumns_block_39__N_1197[5] ), 
         .B(\enc_new_block[19] ), .C(\round_logic.mixcolumns_block_47__N_1397[5] ), 
         .Z(n28939)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i2_3_lut_adj_474.init = 16'h9696;
    LUT4 \round_key_gen.trw_5__bdd_4_lut_29788  (.A(round_key[29]), .B(n11634), 
         .C(n33927), .D(\round_logic.mixcolumns_block_7__N_1245[6] ), .Z(n33091)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam \round_key_gen.trw_5__bdd_4_lut_29788 .init = 16'h6996;
    LUT4 \round_key_gen.trw_5__bdd_3_lut  (.A(\round_key_gen.trw[5] ), .B(n33091), 
         .C(n33846), .Z(n33092)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \round_key_gen.trw_5__bdd_3_lut .init = 16'hcaca;
    LUT4 i1_2_lut_adj_475 (.A(\enc_new_block[57] ), .B(\enc_new_block[17] ), 
         .Z(n11593)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_adj_475.init = 16'h6666;
    PFUMX i28252 (.BLUT(n32321), .ALUT(n32320), .C0(n33847), .Z(n32322));
    PFUMX mux_691_i90 (.BLUT(n2_adj_8034), .ALUT(n5932[89]), .C0(n33843), 
          .Z(n5291[89]));
    LUT4 i27257_3_lut_4_lut (.A(\block_new_127__N_1645[3] ), .B(n33846), 
         .C(n33847), .D(n12936), .Z(n5932[3])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27257_3_lut_4_lut.init = 16'hf808;
    LUT4 i1_2_lut_adj_476 (.A(\round_logic.mixcolumns_block_47__N_1397[6] ), 
         .B(\round_logic.mixcolumns_block_39__N_1197[7] ), .Z(n28869)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_adj_476.init = 16'h6666;
    LUT4 i27255_3_lut_4_lut (.A(\block_new_127__N_1645[2] ), .B(n33846), 
         .C(n33847), .D(n12935), .Z(n5932[2])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27255_3_lut_4_lut.init = 16'hf808;
    LUT4 i1_4_lut_adj_477 (.A(n6347[3]), .B(n33841), .C(n20693), .D(n33847), 
         .Z(block_w1_we)) /* synthesis lut_function=(!(A+!(B (C+(D))+!B !((D)+!C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(422[7] 479[14])
    defparam i1_4_lut_adj_477.init = 16'h4450;
    PFUMX i28240 (.BLUT(n32306), .ALUT(n32305), .C0(n33847), .Z(n32307));
    LUT4 round_key_26__bdd_3_lut (.A(round_key[26]), .B(n33846), .C(\block_reg[3][26] ), 
         .Z(n33108)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_26__bdd_3_lut.init = 16'h4848;
    LUT4 \round_key_gen.trw_2__bdd_4_lut_29807  (.A(round_key[26]), .B(n11630), 
         .C(n11641), .D(\enc_new_block[114] ), .Z(n33110)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam \round_key_gen.trw_2__bdd_4_lut_29807 .init = 16'h6996;
    LUT4 \round_key_gen.trw_2__bdd_3_lut  (.A(\round_key_gen.trw[2] ), .B(n33110), 
         .C(n33846), .Z(n33111)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \round_key_gen.trw_2__bdd_3_lut .init = 16'hcaca;
    LUT4 i1_2_lut_adj_478 (.A(n6347[2]), .B(n6347[3]), .Z(n28866)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_478.init = 16'heeee;
    LUT4 i27253_3_lut_4_lut (.A(\block_new_127__N_1645[1] ), .B(n33846), 
         .C(n33847), .D(n12934), .Z(n5932[1])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27253_3_lut_4_lut.init = 16'hf808;
    LUT4 i20131_2_lut (.A(enc_round_nr[1]), .B(enc_round_nr[0]), .Z(n21[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(387[27:47])
    defparam i20131_2_lut.init = 16'h6666;
    PFUMX i28236 (.BLUT(n32300), .ALUT(n32299), .C0(n33847), .Z(n32301));
    LUT4 i20129_1_lut (.A(enc_round_nr[0]), .Z(n21[0])) /* synthesis lut_function=(!(A)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(387[27:47])
    defparam i20129_1_lut.init = 16'h5555;
    LUT4 round_key_24__bdd_3_lut (.A(round_key[24]), .B(n33846), .C(\block_reg[3][24] ), 
         .Z(n33122)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_24__bdd_3_lut.init = 16'h4848;
    LUT4 \round_key_gen.trw_0__bdd_4_lut_29819  (.A(round_key[24]), .B(n33923), 
         .C(n29080), .D(\enc_new_block[31] ), .Z(n33124)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam \round_key_gen.trw_0__bdd_4_lut_29819 .init = 16'h6996;
    LUT4 \round_key_gen.trw_0__bdd_3_lut  (.A(\round_key_gen.trw[0] ), .B(n33124), 
         .C(n33846), .Z(n33125)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \round_key_gen.trw_0__bdd_3_lut .init = 16'hcaca;
    LUT4 round_key_23__bdd_3_lut (.A(round_key[23]), .B(n33846), .C(\block_reg[3][23] ), 
         .Z(n33131)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_23__bdd_3_lut.init = 16'h4848;
    LUT4 new_sboxw_23__bdd_4_lut (.A(round_key[23]), .B(n28930), .C(\round_logic.mixcolumns_block_15__N_1453[0] ), 
         .D(\enc_new_block[118] ), .Z(n33133)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam new_sboxw_23__bdd_4_lut.init = 16'h6996;
    LUT4 new_sboxw_23__bdd_3_lut (.A(\new_sboxw[23] ), .B(n33133), .C(n33846), 
         .Z(n33134)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam new_sboxw_23__bdd_3_lut.init = 16'hcaca;
    LUT4 i27353_3_lut_4_lut (.A(\block_new_127__N_1645[51] ), .B(n33846), 
         .C(n33847), .D(n12984), .Z(n5932[51])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27353_3_lut_4_lut.init = 16'hf808;
    LUT4 i1_4_lut_adj_479 (.A(n6347[3]), .B(n33841), .C(n20687), .D(n33847), 
         .Z(block_w3_we)) /* synthesis lut_function=(!(A+!(B (C+(D))+!B !((D)+!C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i1_4_lut_adj_479.init = 16'h4450;
    LUT4 i15165_3_lut (.A(n33845), .B(n33846), .C(n6364[3]), .Z(n20687)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i15165_3_lut.init = 16'hdcdc;
    LUT4 round_key_22__bdd_3_lut (.A(round_key[22]), .B(n33846), .C(\block_reg[3][22] ), 
         .Z(n33137)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_22__bdd_3_lut.init = 16'h4848;
    LUT4 new_sboxw_22__bdd_4_lut (.A(round_key[22]), .B(n33928), .C(n33927), 
         .D(\enc_new_block[30] ), .Z(n33139)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam new_sboxw_22__bdd_4_lut.init = 16'h6996;
    LUT4 new_sboxw_22__bdd_3_lut (.A(\new_sboxw[22] ), .B(n33139), .C(n33846), 
         .Z(n33140)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam new_sboxw_22__bdd_3_lut.init = 16'hcaca;
    PFUMX mux_691_i88 (.BLUT(n2_adj_8197), .ALUT(n5932[87]), .C0(n33843), 
          .Z(n5291[87]));
    PFUMX mux_691_i87 (.BLUT(n2_adj_8194), .ALUT(n5932[86]), .C0(n33843), 
          .Z(n5291[86]));
    PFUMX mux_691_i86 (.BLUT(n2_adj_8191), .ALUT(n5932[85]), .C0(n33843), 
          .Z(n5291[85]));
    PFUMX mux_691_i85 (.BLUT(n2_adj_8188), .ALUT(n5932[84]), .C0(n33843), 
          .Z(n5291[84]));
    PFUMX mux_691_i84 (.BLUT(n2_adj_8185), .ALUT(n5932[83]), .C0(n33843), 
          .Z(n5291[83]));
    PFUMX mux_691_i83 (.BLUT(n2_adj_8182), .ALUT(n5932[82]), .C0(n33843), 
          .Z(n5291[82]));
    PFUMX mux_691_i82 (.BLUT(n2_adj_8179), .ALUT(n5932[81]), .C0(n33843), 
          .Z(n5291[81]));
    PFUMX i28230 (.BLUT(n32291), .ALUT(n32290), .C0(n33847), .Z(n32292));
    PFUMX mux_691_i77 (.BLUT(n2_adj_8176), .ALUT(n5932[76]), .C0(n33843), 
          .Z(n5291[76]));
    PFUMX mux_691_i76 (.BLUT(n2_adj_8173), .ALUT(n5932[75]), .C0(n33843), 
          .Z(n5291[75]));
    PFUMX i28226 (.BLUT(n32285), .ALUT(n32284), .C0(n33847), .Z(n32286));
    LUT4 i27351_3_lut_4_lut (.A(\block_new_127__N_1645[50] ), .B(n33846), 
         .C(n33847), .D(n12983), .Z(n5932[50])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27351_3_lut_4_lut.init = 16'hf808;
    PFUMX i28220 (.BLUT(n32276), .ALUT(n32275), .C0(n33847), .Z(n32277));
    PFUMX i28210 (.BLUT(n32262), .ALUT(n32261), .C0(n33847), .Z(n32263));
    PFUMX i28207 (.BLUT(n32256), .ALUT(n32255), .C0(n33847), .Z(n32257));
    PFUMX i28204 (.BLUT(n32250), .ALUT(n32249), .C0(n33847), .Z(n32251));
    PFUMX i28201 (.BLUT(n32244), .ALUT(n32243), .C0(n33847), .Z(n32245));
    PFUMX mux_691_i74 (.BLUT(n2_adj_8170), .ALUT(n5932[73]), .C0(n33843), 
          .Z(n5291[73]));
    PFUMX i28185 (.BLUT(n32224), .ALUT(n32223), .C0(n33847), .Z(n32225));
    PFUMX mux_691_i72 (.BLUT(n2_adj_8167), .ALUT(n5932[71]), .C0(n33843), 
          .Z(n5291[71]));
    LUT4 i27349_3_lut_4_lut (.A(\block_new_127__N_1645[49] ), .B(n33846), 
         .C(n33847), .D(n12982), .Z(n5932[49])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27349_3_lut_4_lut.init = 16'hf808;
    PFUMX mux_691_i71 (.BLUT(n2_adj_8164), .ALUT(n5932[70]), .C0(n33843), 
          .Z(n5291[70]));
    PFUMX mux_691_i70 (.BLUT(n2_adj_8161), .ALUT(n5932[69]), .C0(n33843), 
          .Z(n5291[69]));
    PFUMX mux_691_i69 (.BLUT(n2_adj_8158), .ALUT(n5932[68]), .C0(n33843), 
          .Z(n5291[68]));
    PFUMX i28176 (.BLUT(n32212), .ALUT(n32211), .C0(n33847), .Z(n32213));
    PFUMX mux_691_i68 (.BLUT(n2_adj_8155), .ALUT(n5932[67]), .C0(n33843), 
          .Z(n5291[67]));
    LUT4 round_key_18__bdd_3_lut (.A(round_key[18]), .B(n33846), .C(\block_reg[3][18] ), 
         .Z(n33158)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_18__bdd_3_lut.init = 16'h4848;
    PFUMX mux_691_i66 (.BLUT(n2_adj_8152), .ALUT(n5932[65]), .C0(n33843), 
          .Z(n5291[65]));
    PFUMX mux_691_i65 (.BLUT(n2_adj_8149), .ALUT(n5932[64]), .C0(n33843), 
          .Z(n5291[64]));
    PFUMX i28170 (.BLUT(n32203), .ALUT(n32202), .C0(n33847), .Z(n32204));
    PFUMX mux_691_i63 (.BLUT(n2_adj_8146), .ALUT(n5932[62]), .C0(n33843), 
          .Z(n5291[62]));
    PFUMX mux_691_i62 (.BLUT(n2_adj_8143), .ALUT(n5932[61]), .C0(n33843), 
          .Z(n5291[61]));
    PFUMX mux_691_i61 (.BLUT(n2_adj_8140), .ALUT(n5932[60]), .C0(n33843), 
          .Z(n5291[60]));
    PFUMX mux_691_i60 (.BLUT(n2_adj_8138), .ALUT(n5932[59]), .C0(n33843), 
          .Z(n5291[59]));
    PFUMX mux_691_i58 (.BLUT(n2_adj_8136), .ALUT(n5932[57]), .C0(n33843), 
          .Z(n5291[57]));
    PFUMX i28164 (.BLUT(n32194), .ALUT(n32193), .C0(n33847), .Z(n32195));
    LUT4 new_sboxw_18__bdd_4_lut (.A(round_key[18]), .B(n11641), .C(n33918), 
         .D(\enc_new_block[113] ), .Z(n33160)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam new_sboxw_18__bdd_4_lut.init = 16'h6996;
    LUT4 new_sboxw_18__bdd_3_lut (.A(\new_sboxw[18] ), .B(n33160), .C(n33846), 
         .Z(n33161)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam new_sboxw_18__bdd_3_lut.init = 16'hcaca;
    PFUMX i28157 (.BLUT(n32183), .ALUT(n32182), .C0(n33847), .Z(n32184));
    LUT4 i27339_3_lut_4_lut (.A(\block_new_127__N_1645[44] ), .B(n33846), 
         .C(n33847), .D(n12977), .Z(n5932[44])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27339_3_lut_4_lut.init = 16'hf808;
    LUT4 i27337_3_lut_4_lut (.A(\block_new_127__N_1645[43] ), .B(n33846), 
         .C(n33847), .D(n12976), .Z(n5932[43])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27337_3_lut_4_lut.init = 16'hf808;
    LUT4 i27333_3_lut_4_lut (.A(\block_new_127__N_1645[41] ), .B(n33846), 
         .C(n33847), .D(n12974), .Z(n5932[41])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27333_3_lut_4_lut.init = 16'hf808;
    LUT4 round_key_16__bdd_3_lut (.A(round_key[16]), .B(n33846), .C(\block_reg[3][16] ), 
         .Z(n33172)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_16__bdd_3_lut.init = 16'h4848;
    LUT4 new_sboxw_16__bdd_4_lut (.A(round_key[16]), .B(n33920), .C(n29080), 
         .D(\enc_new_block[24] ), .Z(n33174)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam new_sboxw_16__bdd_4_lut.init = 16'h6996;
    LUT4 new_sboxw_16__bdd_3_lut (.A(\new_sboxw[16] ), .B(n33174), .C(n33846), 
         .Z(n33175)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam new_sboxw_16__bdd_3_lut.init = 16'hcaca;
    LUT4 round_key_15__bdd_3_lut (.A(round_key[15]), .B(n33846), .C(\block_reg[3][15] ), 
         .Z(n33181)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_15__bdd_3_lut.init = 16'h4848;
    LUT4 i27329_3_lut_4_lut (.A(\block_new_127__N_1645[39] ), .B(n33846), 
         .C(n33847), .D(n12972), .Z(n5932[39])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27329_3_lut_4_lut.init = 16'hf808;
    PFUMX i28154 (.BLUT(n32177), .ALUT(n32176), .C0(n33847), .Z(n32178));
    LUT4 i27325_3_lut_4_lut (.A(\block_new_127__N_1645[37] ), .B(n33846), 
         .C(n33847), .D(n12970), .Z(n5932[37])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27325_3_lut_4_lut.init = 16'hf808;
    LUT4 i27323_3_lut_4_lut (.A(\block_new_127__N_1645[36] ), .B(n33846), 
         .C(n33847), .D(n12969), .Z(n5932[36])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27323_3_lut_4_lut.init = 16'hf808;
    LUT4 \round_key_gen.trw_23__bdd_4_lut_29685  (.A(round_key[15]), .B(n28930), 
         .C(\enc_new_block[119] ), .D(\round_logic.mixcolumns_block_7__N_1245[7] ), 
         .Z(n33183)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam \round_key_gen.trw_23__bdd_4_lut_29685 .init = 16'h6996;
    LUT4 \round_key_gen.trw_23__bdd_3_lut  (.A(\round_key_gen.trw[23] ), .B(n33183), 
         .C(n33846), .Z(n33184)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \round_key_gen.trw_23__bdd_3_lut .init = 16'hcaca;
    PFUMX mux_691_i52 (.BLUT(n2_adj_8133), .ALUT(n5932[51]), .C0(n33843), 
          .Z(n5291[51]));
    PFUMX mux_691_i51 (.BLUT(n2_adj_8130), .ALUT(n5932[50]), .C0(n33843), 
          .Z(n5291[50]));
    LUT4 i27319_3_lut_4_lut (.A(\block_new_127__N_1645[34] ), .B(n33846), 
         .C(n33847), .D(n12967), .Z(n5932[34])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27319_3_lut_4_lut.init = 16'hf808;
    LUT4 round_key_13__bdd_3_lut (.A(round_key[13]), .B(n33846), .C(\block_reg[3][13] ), 
         .Z(n33193)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_13__bdd_3_lut.init = 16'h4848;
    PFUMX mux_691_i50 (.BLUT(n2_adj_8127), .ALUT(n5932[49]), .C0(n33843), 
          .Z(n5291[49]));
    LUT4 i27317_3_lut_4_lut (.A(\block_new_127__N_1645[33] ), .B(n33846), 
         .C(n33847), .D(n12966), .Z(n5932[33])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27317_3_lut_4_lut.init = 16'hf808;
    LUT4 \round_key_gen.trw_21__bdd_4_lut_29696  (.A(round_key[13]), .B(n33921), 
         .C(n33919), .D(\enc_new_block[117] ), .Z(n33195)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam \round_key_gen.trw_21__bdd_4_lut_29696 .init = 16'h6996;
    LUT4 \round_key_gen.trw_21__bdd_3_lut  (.A(\round_key_gen.trw[21] ), .B(n33195), 
         .C(n33846), .Z(n33196)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \round_key_gen.trw_21__bdd_3_lut .init = 16'hcaca;
    LUT4 i27311_3_lut_4_lut (.A(\block_new_127__N_1645[30] ), .B(n33846), 
         .C(n33847), .D(n12963), .Z(n5932[30])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27311_3_lut_4_lut.init = 16'hf808;
    LUT4 round_key_11__bdd_3_lut (.A(round_key[11]), .B(n33846), .C(\block_reg[3][11] ), 
         .Z(n33205)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_11__bdd_3_lut.init = 16'h4848;
    LUT4 i27307_3_lut_4_lut (.A(\block_new_127__N_1645[28] ), .B(n33846), 
         .C(n33847), .D(n12961), .Z(n5932[28])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27307_3_lut_4_lut.init = 16'hf808;
    LUT4 i27305_3_lut_4_lut (.A(\block_new_127__N_1645[27] ), .B(n33846), 
         .C(n33847), .D(n12960), .Z(n5932[27])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27305_3_lut_4_lut.init = 16'hf808;
    LUT4 \round_key_gen.trw_19__bdd_3_lut  (.A(\round_key_gen.trw[19] ), .B(n33207), 
         .C(n33846), .Z(n33208)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \round_key_gen.trw_19__bdd_3_lut .init = 16'hcaca;
    LUT4 i1_4_lut_adj_480 (.A(n6347[3]), .B(n33841), .C(n20696), .D(n33847), 
         .Z(block_w0_we)) /* synthesis lut_function=(!(A+!(B (C+(D))+!B !((D)+!C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(422[7] 479[14])
    defparam i1_4_lut_adj_480.init = 16'h4450;
    LUT4 round_key_9__bdd_3_lut (.A(round_key[9]), .B(n33846), .C(\block_reg[3][9] ), 
         .Z(n33217)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_9__bdd_3_lut.init = 16'h4848;
    LUT4 i15174_3_lut (.A(n33845), .B(n33846), .C(n6364_c[0]), .Z(n20696)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i15174_3_lut.init = 16'hdcdc;
    LUT4 i27301_3_lut_4_lut (.A(\block_new_127__N_1645[25] ), .B(n33846), 
         .C(n33847), .D(n12958), .Z(n5932[25])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27301_3_lut_4_lut.init = 16'hf808;
    PFUMX mux_691_i45 (.BLUT(n2_adj_8122), .ALUT(n5932[44]), .C0(n33843), 
          .Z(n5291[44]));
    LUT4 \round_key_gen.trw_17__bdd_4_lut_29720  (.A(round_key[9]), .B(n33853), 
         .C(n11630), .D(n33917), .Z(n33219)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam \round_key_gen.trw_17__bdd_4_lut_29720 .init = 16'h6996;
    LUT4 \round_key_gen.trw_17__bdd_3_lut  (.A(\round_key_gen.trw[17] ), .B(n33219), 
         .C(n33846), .Z(n33220)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \round_key_gen.trw_17__bdd_3_lut .init = 16'hcaca;
    LUT4 round_key_8__bdd_3_lut (.A(round_key[8]), .B(n33846), .C(\block_reg[3][8] ), 
         .Z(n33223)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_8__bdd_3_lut.init = 16'h4848;
    LUT4 \round_key_gen.trw_16__bdd_3_lut  (.A(\round_key_gen.trw[16] ), .B(n33225), 
         .C(n33846), .Z(n33226)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \round_key_gen.trw_16__bdd_3_lut .init = 16'hcaca;
    PFUMX mux_691_i44 (.BLUT(n2_adj_8119), .ALUT(n5932[43]), .C0(n33843), 
          .Z(n5291[43]));
    PFUMX mux_691_i42 (.BLUT(n2_adj_8107), .ALUT(n5932[41]), .C0(n33843), 
          .Z(n5291[41]));
    PFUMX mux_691_i40 (.BLUT(n2_adj_8098), .ALUT(n5932[39]), .C0(n33843), 
          .Z(n5291[39]));
    LUT4 round_key_6__bdd_3_lut (.A(round_key[6]), .B(n33846), .C(\block_reg[3][6] ), 
         .Z(n33235)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_6__bdd_3_lut.init = 16'h4848;
    LUT4 i27293_3_lut_4_lut (.A(\block_new_127__N_1645[21] ), .B(n33846), 
         .C(n33847), .D(n12954), .Z(n5932[21])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27293_3_lut_4_lut.init = 16'hf808;
    LUT4 \round_key_gen.trw_14__bdd_4_lut_29746  (.A(round_key[6]), .B(n33930), 
         .C(n33921), .D(\round_logic.mixcolumns_block_15__N_1453[7] ), .Z(n33237)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam \round_key_gen.trw_14__bdd_4_lut_29746 .init = 16'h6996;
    LUT4 \round_key_gen.trw_14__bdd_3_lut  (.A(\round_key_gen.trw[14] ), .B(n33237), 
         .C(n33846), .Z(n33238)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \round_key_gen.trw_14__bdd_3_lut .init = 16'hcaca;
    PFUMX mux_691_i38 (.BLUT(n2_adj_8083), .ALUT(n5932[37]), .C0(n33843), 
          .Z(n5291[37]));
    LUT4 i27291_3_lut_4_lut (.A(\block_new_127__N_1645[20] ), .B(n33846), 
         .C(n33847), .D(n12953), .Z(n5932[20])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27291_3_lut_4_lut.init = 16'hf808;
    LUT4 i27289_3_lut_4_lut (.A(\block_new_127__N_1645[19] ), .B(n33846), 
         .C(n33847), .D(n12952), .Z(n5932[19])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27289_3_lut_4_lut.init = 16'hf808;
    LUT4 i27285_3_lut_4_lut (.A(\block_new_127__N_1645[17] ), .B(n33846), 
         .C(n33847), .D(n12950), .Z(n5932[17])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27285_3_lut_4_lut.init = 16'hf808;
    PFUMX mux_691_i37 (.BLUT(n2_adj_8064), .ALUT(n5932[36]), .C0(n33843), 
          .Z(n5291[36]));
    PFUMX mux_691_i35 (.BLUT(n2_adj_8055), .ALUT(n5932[34]), .C0(n33843), 
          .Z(n5291[34]));
    PFUMX mux_691_i34 (.BLUT(n2_adj_8052), .ALUT(n5932[33]), .C0(n33843), 
          .Z(n5291[33]));
    PFUMX mux_691_i31 (.BLUT(n2_adj_8049), .ALUT(n5932[30]), .C0(n33843), 
          .Z(n5291[30]));
    PFUMX mux_691_i29 (.BLUT(n2_adj_8046), .ALUT(n5932[28]), .C0(n33843), 
          .Z(n5291[28]));
    PFUMX mux_691_i28 (.BLUT(n2_adj_8043), .ALUT(n5932[27]), .C0(n33843), 
          .Z(n5291[27]));
    LUT4 i27279_3_lut_4_lut (.A(\block_new_127__N_1645[14] ), .B(n33846), 
         .C(n33847), .D(n12947), .Z(n5932[14])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(281[7] 343[14])
    defparam i27279_3_lut_4_lut.init = 16'hf808;
    PFUMX mux_691_i26 (.BLUT(n2_adj_8031), .ALUT(n5932[25]), .C0(n33843), 
          .Z(n5291[25]));
    LUT4 round_key_0__bdd_3_lut (.A(round_key[0]), .B(n33846), .C(\block_reg[3][0] ), 
         .Z(n33270)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam round_key_0__bdd_3_lut.init = 16'h4848;
    LUT4 \round_key_gen.trw_8__bdd_4_lut_29775  (.A(round_key[0]), .B(n33922), 
         .C(n12156), .D(\enc_new_block[72] ), .Z(n33272)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam \round_key_gen.trw_8__bdd_4_lut_29775 .init = 16'h6996;
    LUT4 \round_key_gen.trw_8__bdd_3_lut  (.A(\round_key_gen.trw[8] ), .B(n33272), 
         .C(n33846), .Z(n33273)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \round_key_gen.trw_8__bdd_3_lut .init = 16'hcaca;
    PFUMX mux_691_i22 (.BLUT(n2_adj_8030), .ALUT(n5932[21]), .C0(n33843), 
          .Z(n5291[21]));
    PFUMX mux_691_i21 (.BLUT(n2_adj_8027), .ALUT(n5932[20]), .C0(n33843), 
          .Z(n5291[20]));
    LUT4 i1_2_lut_adj_481 (.A(\enc_new_block[87] ), .B(\round_logic.mixcolumns_block_103__N_1101[0] ), 
         .Z(n29399)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_adj_481.init = 16'h6666;
    LUT4 i2_2_lut_adj_482 (.A(\round_logic.mixcolumns_block_103__N_1101[6] ), 
         .B(\enc_new_block[84] ), .Z(n7_adj_8114)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i2_2_lut_adj_482.init = 16'h6666;
    PFUMX mux_691_i20 (.BLUT(n2), .ALUT(n5932[19]), .C0(n33843), .Z(n5291[19]));
    LUT4 i3_3_lut_adj_483 (.A(n29105), .B(\enc_new_block[122] ), .C(round_key[123]), 
         .Z(n8_adj_8112)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i3_3_lut_adj_483.init = 16'h9696;
    LUT4 i2_3_lut_adj_484 (.A(\enc_new_block[43] ), .B(\enc_new_block[82] ), 
         .C(\enc_new_block[3] ), .Z(n29105)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i2_3_lut_adj_484.init = 16'h9696;
    LUT4 i2_2_lut_adj_485 (.A(round_key[121]), .B(\enc_new_block[81] ), 
         .Z(n7_adj_8108)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(87[13:53])
    defparam i2_2_lut_adj_485.init = 16'h6666;
    LUT4 i1_2_lut_adj_486 (.A(\enc_new_block[40] ), .B(\enc_new_block[80] ), 
         .Z(n29077)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i1_2_lut_adj_486.init = 16'h6666;
    PFUMX mux_691_i18 (.BLUT(n2_adj_8228), .ALUT(n5932[17]), .C0(n33843), 
          .Z(n5291[17]));
    PFUMX mux_691_i15 (.BLUT(n2_adj_8226), .ALUT(n5932[14]), .C0(n33843), 
          .Z(n5291[14]));
    PFUMX mux_691_i13 (.BLUT(n2_adj_8224), .ALUT(n5932[12]), .C0(n33843), 
          .Z(n5291[12]));
    LUT4 i2_2_lut_adj_487 (.A(\round_logic.mixcolumns_block_111__N_1285[7] ), 
         .B(\round_logic.mixcolumns_block_111__N_1285[0] ), .Z(n7_adj_8102)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(153[21:32])
    defparam i2_2_lut_adj_487.init = 16'h6666;
    PFUMX mux_691_i11 (.BLUT(n2_adj_8221), .ALUT(n5932[10]), .C0(n33843), 
          .Z(n5291[10]));
    PFUMX mux_691_i8 (.BLUT(n2_adj_8219), .ALUT(n5932[7]), .C0(n33843), 
          .Z(n5291[7]));
    PFUMX mux_691_i6 (.BLUT(n2_adj_8217), .ALUT(n5932[5]), .C0(n33843), 
          .Z(n5291[5]));
    PFUMX mux_691_i5 (.BLUT(n2_adj_8215), .ALUT(n5932[4]), .C0(n33843), 
          .Z(n5291[4]));
    PFUMX mux_691_i4 (.BLUT(n2_adj_8213), .ALUT(n5932[3]), .C0(n33843), 
          .Z(n5291[3]));
    PFUMX mux_691_i3 (.BLUT(n2_adj_8211), .ALUT(n5932[2]), .C0(n33843), 
          .Z(n5291[2]));
    PFUMX mux_691_i2 (.BLUT(n2_adj_8209), .ALUT(n5932[1]), .C0(n33843), 
          .Z(n5291[1]));
    
endmodule
//
// Verilog Description of module aes_decipher_block
//

module aes_decipher_block (dec_new_block, round_key, clk_c, tmp_sboxw, 
            dec_round_nr, round_ctr_we, round_ctr_new, n6347, encdec_reg, 
            \aes_core_ctrl_new_1__N_858[1] , n28773, \enc_round_nr[3] , 
            block_w3_we_N_1490, n4, n33858, n149, block_new_127__N_1645, 
            \block_new_127__N_1645[37] , \block_new_127__N_1645[36] , \block_new_127__N_1645[34] , 
            \block_new_127__N_1645[33] , \block_new_127__N_1645[62] , \block_new_127__N_1645[61] , 
            \block_new_127__N_1645[60] , \block_new_127__N_1645[59] , \block_new_127__N_1645[57] , 
            \block_new_127__N_1645[87] , \block_new_127__N_1645[86] , \block_new_127__N_1645[85] , 
            \block_new_127__N_1645[84] , \block_new_127__N_1645[83] , \block_new_127__N_1645[82] , 
            \block_new_127__N_1645[81] , \block_new_127__N_1645[108] , \block_new_127__N_1645[107] , 
            \block_new_127__N_1645[105] , \block_new_127__N_1645[7] , \block_new_127__N_1645[5] , 
            \block_new_127__N_1645[4] , \block_new_127__N_1645[3] , \block_new_127__N_1645[2] , 
            \enc_round_nr[1] , \muxed_round_nr[1] , \block_new_127__N_1645[1] , 
            \block_new_127__N_1645[30] , new_sboxw, \block_new_127__N_1645[28] , 
            \block_new_127__N_1645[27] , \block_new_127__N_1645[25] , \block_reg[0] , 
            \block_new_127__N_1645[51] , \block_new_127__N_1645[50] , \block_new_127__N_1645[49] , 
            dec_ready, dec_ctrl_we, \block_new_127__N_1645[76] , \block_new_127__N_1645[125] , 
            \block_new_127__N_1645[123] , \key_mem_ctrl.num_rounds[2] , 
            \muxed_round_nr[3] , \enc_round_nr[2] , \muxed_round_nr[2] , 
            \block_new_127__N_1645[121] , \block_new_127__N_1645[21] , \block_new_127__N_1645[20] , 
            \block_new_127__N_1645[19] , \block_new_127__N_1645[17] , \block_new_127__N_1645[44] , 
            \block_new_127__N_1645[43] , \block_new_127__N_1645[41] , \block_new_127__N_1645[71] , 
            \block_new_127__N_1645[70] , \block_new_127__N_1645[69] , \block_new_127__N_1645[68] , 
            \block_new_127__N_1645[67] , \block_new_127__N_1645[65] , \block_new_127__N_1645[64] , 
            \block_new_127__N_1645[92] , \block_new_127__N_1645[91] , \block_new_127__N_1645[89] , 
            \block_new_127__N_1645[119] , \block_new_127__N_1645[118] , 
            \block_new_127__N_1645[116] , \block_new_127__N_1645[115] , 
            \block_new_127__N_1645[114] , \block_new_127__N_1645[113] , 
            \block_new_127__N_1645[14] , \block_new_127__N_1645[12] , \block_new_127__N_1645[10] , 
            \block_new_127__N_1645[75] , \block_new_127__N_1645[73] , \block_new_127__N_1645[102] , 
            \block_new_127__N_1645[99] , \block_new_127__N_1645[98] , \block_new_127__N_1645[97] , 
            n14934, dec_ctrl_new_2__N_2032, n33848, n33846, \block_reg[1] , 
            \block_reg[3] , \round_ctr_new[3] , n33942, n33913, enc_ready, 
            n6428, \block_reg[2] , n14930, n33909, n14939, n152) /* synthesis syn_module_defined=1 */ ;
    output [127:0]dec_new_block;
    input [127:0]round_key;
    input clk_c;
    output [31:0]tmp_sboxw;
    output [3:0]dec_round_nr;
    input round_ctr_we;
    input [3:0]round_ctr_new;
    input [3:0]n6347;
    input encdec_reg;
    input \aes_core_ctrl_new_1__N_858[1] ;
    output n28773;
    input \enc_round_nr[3] ;
    input block_w3_we_N_1490;
    input n4;
    input n33858;
    output n149;
    output [127:0]block_new_127__N_1645;
    output \block_new_127__N_1645[37] ;
    output \block_new_127__N_1645[36] ;
    output \block_new_127__N_1645[34] ;
    output \block_new_127__N_1645[33] ;
    output \block_new_127__N_1645[62] ;
    output \block_new_127__N_1645[61] ;
    output \block_new_127__N_1645[60] ;
    output \block_new_127__N_1645[59] ;
    output \block_new_127__N_1645[57] ;
    output \block_new_127__N_1645[87] ;
    output \block_new_127__N_1645[86] ;
    output \block_new_127__N_1645[85] ;
    output \block_new_127__N_1645[84] ;
    output \block_new_127__N_1645[83] ;
    output \block_new_127__N_1645[82] ;
    output \block_new_127__N_1645[81] ;
    output \block_new_127__N_1645[108] ;
    output \block_new_127__N_1645[107] ;
    output \block_new_127__N_1645[105] ;
    output \block_new_127__N_1645[7] ;
    output \block_new_127__N_1645[5] ;
    output \block_new_127__N_1645[4] ;
    output \block_new_127__N_1645[3] ;
    output \block_new_127__N_1645[2] ;
    input \enc_round_nr[1] ;
    output \muxed_round_nr[1] ;
    output \block_new_127__N_1645[1] ;
    output \block_new_127__N_1645[30] ;
    input [31:0]new_sboxw;
    output \block_new_127__N_1645[28] ;
    output \block_new_127__N_1645[27] ;
    output \block_new_127__N_1645[25] ;
    input [31:0]\block_reg[0] ;
    output \block_new_127__N_1645[51] ;
    output \block_new_127__N_1645[50] ;
    output \block_new_127__N_1645[49] ;
    output dec_ready;
    input dec_ctrl_we;
    output \block_new_127__N_1645[76] ;
    output \block_new_127__N_1645[125] ;
    output \block_new_127__N_1645[123] ;
    input \key_mem_ctrl.num_rounds[2] ;
    output \muxed_round_nr[3] ;
    input \enc_round_nr[2] ;
    output \muxed_round_nr[2] ;
    output \block_new_127__N_1645[121] ;
    output \block_new_127__N_1645[21] ;
    output \block_new_127__N_1645[20] ;
    output \block_new_127__N_1645[19] ;
    output \block_new_127__N_1645[17] ;
    output \block_new_127__N_1645[44] ;
    output \block_new_127__N_1645[43] ;
    output \block_new_127__N_1645[41] ;
    output \block_new_127__N_1645[71] ;
    output \block_new_127__N_1645[70] ;
    output \block_new_127__N_1645[69] ;
    output \block_new_127__N_1645[68] ;
    output \block_new_127__N_1645[67] ;
    output \block_new_127__N_1645[65] ;
    output \block_new_127__N_1645[64] ;
    output \block_new_127__N_1645[92] ;
    output \block_new_127__N_1645[91] ;
    output \block_new_127__N_1645[89] ;
    output \block_new_127__N_1645[119] ;
    output \block_new_127__N_1645[118] ;
    output \block_new_127__N_1645[116] ;
    output \block_new_127__N_1645[115] ;
    output \block_new_127__N_1645[114] ;
    output \block_new_127__N_1645[113] ;
    output \block_new_127__N_1645[14] ;
    output \block_new_127__N_1645[12] ;
    output \block_new_127__N_1645[10] ;
    output \block_new_127__N_1645[75] ;
    output \block_new_127__N_1645[73] ;
    output \block_new_127__N_1645[102] ;
    output \block_new_127__N_1645[99] ;
    output \block_new_127__N_1645[98] ;
    output \block_new_127__N_1645[97] ;
    input n14934;
    output dec_ctrl_new_2__N_2032;
    input n33848;
    output n33846;
    input [31:0]\block_reg[1] ;
    input [31:0]\block_reg[3] ;
    input \round_ctr_new[3] ;
    input n33942;
    input n33913;
    input enc_ready;
    output n6428;
    input [31:0]\block_reg[2] ;
    output n14930;
    output n33909;
    output n14939;
    output n152;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(41[33:36])
    
    wire n33756, block_w3_we;
    wire [127:0]n3899;
    wire [31:0]n2752;
    
    wire n9418, n30146, n25333, n33704;
    wire [127:0]block_new_127__N_1901;
    
    wire n5, n33755, n33754, n33753, n33752, n29254, n29172, n29483, 
        n6, n33751, n33750, n33749, n33748, n28961, n33524, n28926, 
        n33506, n12084, n29447, n33523, n33507, n33522, block_w1_we, 
        block_w0_we, n9416, n4_c, n33829;
    wire [7:0]n6228;
    
    wire n33508, n33673, n33686, n33825, n8;
    wire [3:0]dec_round_nr_c;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(99[18:30])
    wire [3:0]round_ctr_new_c;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(201[17:30])
    wire [2:0]update_type;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(230[17:28])
    
    wire n33844, n13131;
    wire [127:0]n4540;
    wire [127:0]block_new_127__N_1645_c;
    
    wire n13130, n13129, n13128, n13127, n13126, n13125, n13124, 
        n13123, n33774, n9, n13122, n13121, n33679, n33766, n33768, 
        n4_adj_7671, n13120, n9394, n33675;
    wire [7:0]n4770;
    
    wire n4_adj_7672, n13119, n13118, n9392, n9_adj_7673, n13117, 
        n13116, n9414, n9390, n7, n13115, n29441, n8_adj_7674;
    wire [7:0]n873;
    wire [7:0]n648;
    
    wire n33509, n9388, n33796, n33803, n9_adj_7675, n13114, n9386, 
        n13113, n13112, n9384, n9382, n8_adj_7676, n9380, n33678, 
        n33688, n7_adj_7677, n33804, n33681, n7_adj_7678, n33692, 
        n33702, n6_adj_7679, n9412, n13111, n13110, n33820, n4_adj_7680, 
        n9378, n13109, n5_adj_7681, n13108, n13107, n13106, n9376, 
        n13105, n33683, n33703, n29381, n8_adj_7682, n33785, n33794, 
        n6_adj_7683, n9374, n13104, n9372, n13103, n13102, n9370, 
        n33699, n33706, n33684, n8_adj_7684, n13101, n13100, n13099, 
        n13098, n9368, n13097, n33801, n33772, n6_adj_7685, n13096, 
        n13095, n33707, n8_adj_7686, n13094, n33689, n8_adj_7687, 
        n33836, n29160, n33838, n8_adj_7688, n13093, n13092, n9366, 
        n8522, n33763, n33800, n33685, n6_adj_7689, n33786, n11, 
        n28987, n4_adj_7690, n6_adj_7691, n33813, n5_adj_7692, n13091, 
        n33791, n6_adj_7693, n13090, n9410, n8_adj_7694, n5_adj_7695, 
        n2, n5_adj_7696, n6_adj_7697, n2_adj_7698, n4_adj_7699, n7_adj_7700, 
        n8_adj_7701, n2_adj_7702, n6_adj_7703, n2_adj_7704, n29390, 
        n2_adj_7705, n2_adj_7706, n9_adj_7707, n10, n2_adj_7708, n33518, 
        n7_adj_7709, n2_adj_7710, n10_adj_7711, n2_adj_7712, n5_adj_7713, 
        n6_adj_7714, n2_adj_7715, n7_adj_7716, n2_adj_7717, n33690, 
        n33589, n8_adj_7718, n5_adj_7719, n6_adj_7720, n2_adj_7721, 
        n29396, n4_adj_7722, n2_adj_7723, n7_adj_7724, n8_adj_7725, 
        n2_adj_7726, n7_adj_7727, n8_adj_7728, n2_adj_7729, n33781, 
        n33757, n7_adj_7730, n13089, n13088, n33710, n33839, n8_adj_7731, 
        n7_adj_7732, n8_adj_7733, n2_adj_7734, n9_adj_7735, n10_adj_7736, 
        n2_adj_7737, n13087, n33582, n4_adj_7738, n2_adj_7739, n13086, 
        n10_adj_7740, n2_adj_7741, n13085, n5_adj_7742, n6_adj_7743, 
        n2_adj_7744, n9_adj_7745, n10_adj_7746, n2_adj_7747, n33580, 
        n4_adj_7748, n2_adj_7749, n13084, n29375, n4_adj_7750, n2_adj_7751, 
        n5_adj_7752;
    wire [3:0]n6362;
    
    wire n7_adj_7753, n8_adj_7754, n2_adj_7755, n13083, n13082, n7_adj_7756, 
        n2_adj_7757, n33668, n8_adj_7758, n10_adj_7759, n2_adj_7760, 
        n5_adj_7761, n6_adj_7762, n2_adj_7763, n33677, n12090, n13081, 
        n8_adj_7764, n2_adj_7765, n13080, n13079, n4_adj_7766, n2_adj_7767, 
        n13078, n33713, n6_adj_7768, n9408;
    wire [7:0]n3564;
    
    wire n5_adj_7769, n2_adj_7770, n5_adj_7771, n2_adj_7772, n12, 
        n2_adj_7773, n5_adj_7774, n6_adj_7775, n2_adj_7776, n13077, 
        n5_adj_7777, n6_adj_7778, n2_adj_7779, n5_adj_7780, n2_adj_7781, 
        block_w2_we, n9406, n33672, n7_adj_7782, n2_adj_7783, n13076, 
        n29429, n2_adj_7784, n5_adj_7785, n6_adj_7786, n2_adj_7787, 
        n7_adj_7788, n8_adj_7789, n2_adj_7790, n9_adj_7791, n10_adj_7792, 
        n2_adj_7793, sword_ctr_we;
    wire [3:0]n2689;
    
    wire n7_adj_7794, n8_adj_7795, n2_adj_7796, n6_adj_7797, n2_adj_7798, 
        n33583, n33579, n13075, n5_adj_7799, n6_adj_7800, n2_adj_7801, 
        n9396, n9398, n33697, n33587, n33779, n8_adj_7802, n5_adj_7803, 
        n6_adj_7804, n2_adj_7805, n9404, n9400, n5_adj_7806, n6_adj_7807, 
        n2_adj_7808, n5_adj_7809, n6_adj_7810, n2_adj_7811, n33584, 
        n7_adj_7812, n33762, n4_adj_7813, n29273, n4_adj_7814, n2_adj_7815, 
        n9402, n6_adj_7816, n9_adj_7817, n10_adj_7818, n2_adj_7819, 
        n33828, n4_adj_7820, n33698, n33671, n5_adj_7821, n6_adj_7822, 
        n2_adj_7823, n8_adj_7824, n2_adj_7825, n33769, n4_adj_7826, 
        n2_adj_7827, n33520, n2_adj_7828, n33586, n33812, n33799, 
        n8_adj_7829, n9_adj_7830, n10_adj_7831, n2_adj_7832, n6431, 
        n9_adj_7833, n10_adj_7834, n2_adj_7835, n5_adj_7836, n6_adj_7837, 
        n2_adj_7838, n28882, n4_adj_7839, n2_adj_7840, n33519, n4_adj_7841, 
        n2_adj_7842, n4_adj_7843;
    wire [3:0]n6363;
    
    wire n5_adj_7844, n6_adj_7845, n2_adj_7846, n7_adj_7847, n8_adj_7848, 
        n2_adj_7849, n7_adj_7850, n8_adj_7851, n2_adj_7852, n5_adj_7853, 
        n6_adj_7854, n2_adj_7855, n9420, n5_adj_7856, n2_adj_7857, 
        n13074, n29244, n4_adj_7858, n2_adj_7859, n9422, n7_adj_7860, 
        n2_adj_7861, n13187, n7_adj_7862, n2_adj_7863, n13186, n9424, 
        n5_adj_7864, n2_adj_7865, n9_adj_7866, n10_adj_7867, n2_adj_7868, 
        n9426, n13073, n13072, n29291, n4_adj_7869, n2_adj_7870, 
        n33590, n7_adj_7871, n4_adj_7872, n2_adj_7873, n13185, n13184, 
        n7_adj_7874, n8_adj_7875, n2_adj_7876, n14912, n13183, n7_adj_7877, 
        n8_adj_7878, n2_adj_7879, n30080, n110, n13182, n13181, 
        n13180, n7_adj_7880, n8_adj_7881, n2_adj_7882, n7_adj_7883, 
        n2_adj_7884, n5_adj_7885, n6_adj_7886, n2_adj_7887, n13179, 
        n7_adj_7888, n8_adj_7889, n2_adj_7890, n13178, n13177, n29462, 
        n4_adj_7891, n2_adj_7892, n33521, n4_adj_7893, n2_adj_7894, 
        n13176, n13175, n13174, n13173, n13172, n13171, n13170, 
        n13169, n13168, n13167, n13166, n13165, n13164, n13163, 
        n13162, n13161, n13160, n13159, n13158, n13157, n13156, 
        n13155, n13154, n13153, n13152, n13151, n13150, n13149, 
        n13148, n13147, n13146, n13145, n13144, n13143, n13142, 
        n13141, n13140, n13139, n13138, n13137, n13136, n33674, 
        n33782, n13135, n13134, n13133, n33758, n13132, n5_adj_7896, 
        n6_adj_7897, n2_adj_7898, n33693, n4_adj_7899, n2_adj_7900, 
        n5_adj_7901, n6_adj_7902, n2_adj_7903, n33773, n2_adj_7904, 
        n33777, n4_adj_7905, n2_adj_7906, n29444, n33808, n5_adj_7907, 
        n5_adj_7908, n6_adj_7909, n2_adj_7910, n33807, n7_adj_7911, 
        n2_adj_7912, n8_adj_7913, n2_adj_7914, n5_adj_7915, n6_adj_7916, 
        n2_adj_7917, n5_adj_7918, n6_adj_7919, n2_adj_7920, n4_adj_7921, 
        n2_adj_7922, n33790, n33715, n33701, n33837, n6_adj_7923, 
        n5_adj_7924, n2_adj_7925, n5_adj_7926, n6_adj_7927, n2_adj_7928, 
        n6_adj_7929, n2_adj_7930, n33585, n2_adj_7931, n4_adj_7932, 
        n2_adj_7933, n7_adj_7934, n2_adj_7935, n5_adj_7936, n6_adj_7937, 
        n2_adj_7938, n6_adj_7939, n2_adj_7940, n13071, n6_adj_7941, 
        n2_adj_7942, n7_adj_7943, n8_adj_7944, n2_adj_7945, n5_adj_7946, 
        n6_adj_7947, n2_adj_7948, n7_adj_7949, n8_adj_7950, n2_adj_7951, 
        n13070, n5_adj_7952, n6_adj_7953, n2_adj_7954, n33792, n33793, 
        n5_adj_7955, n6_adj_7956, n2_adj_7957, n12748, n7_adj_7958, 
        n33705, n13069, n13068, n13067, n33797, n33588, n13066, 
        n13065, n13064, n33525, n4_adj_7959, n2_adj_7960, n4_adj_7961, 
        n2_adj_7962, n8_adj_7963, n2_adj_7964, n5_adj_7965, n6_adj_7966, 
        n2_adj_7967, n7_adj_7968, n8_adj_7969, n2_adj_7970, n4_adj_7971, 
        n2_adj_7972, n7_adj_7973, n2_adj_7974, n7_adj_7975, n8_adj_7976, 
        n2_adj_7977, n29339, n5_adj_7978, n6_adj_7979, n2_adj_7980, 
        n13063, n13062, n33708, n13061, n33767, n14933, n33676, 
        n29143, n33682, n33669, n33784, n33842, n20699, n29393, 
        n33826, n5_adj_7981, n5_adj_7982, n2_adj_7983, n7_adj_7984, 
        n8_adj_7985, n2_adj_7986, n9_adj_7987, n10_adj_7988, n2_adj_7989, 
        n33780, n5_adj_7990, n2_adj_7991, n7_adj_7992, n2_adj_7993, 
        n5_adj_7994, n2_adj_7995, n33830, n7_adj_7996, n2_adj_7997, 
        n33849, n33935, n20702, n20708, n20705, n33760, n4_adj_7998, 
        n33714, n33691, n33695, n33776, n6_adj_7999, n12810, n12933, 
        n33783, n29288, n33700, n33798, n33687, n11918, n33788, 
        n33823, n33817, n33761, n33574, n33856, n33578, n33806;
    wire [7:0]n5085;
    
    wire n33575;
    wire [7:0]n6327;
    
    wire n8_adj_8000, n33831, n8_adj_8001, n33581, n33809, n33822, 
        n33764, n10_adj_8002, n12_adj_8003, n33795, n33680, n33821, 
        n33816, n33577, n33840, n33576, n2_adj_8004, n14890, n33835, 
        n12921, n33670, n33814, n33805, n29408, n7_adj_8005, n33711, 
        n12071, n2_adj_8006, n33834, n33833, n2_adj_8007, n33832, 
        n29146, n33787, n6_adj_8008, n2_adj_8009, n9_adj_8010, n2_adj_8011, 
        n6_adj_8012, n2_adj_8013, n33827, n33824, n2_adj_8014, n2_adj_8015, 
        n12074, n33819, n33818, n2_adj_8016, n29480, n33694, n11_adj_8017, 
        n33709, n33815, n33811, n33810, n14919, n11890, n33802, 
        n2886, n33789, n33778, n33775, n33771, n33770, n33765, 
        n33759, n28836, n30026, n33936, n29231, n33712, n29471, 
        n6_adj_8018, n166, n2_adj_8019, n6_adj_8020, n29220;
    wire [7:0]n6111;
    
    wire n9_adj_8021, n8_adj_8022;
    wire [7:0]n6345;
    
    wire n29181, n29199, n29432, n6_adj_8023;
    wire [7:0]n6048;
    
    wire n12_adj_8024;
    
    LUT4 i1_2_lut_rep_452_4_lut (.A(dec_new_block[96]), .B(round_key[96]), 
         .C(dec_new_block[112]), .D(round_key[112]), .Z(n33756)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_rep_452_4_lut.init = 16'h6996;
    FD1P3AX block_w3_reg__i1 (.D(n3899[0]), .SP(block_w3_we), .CK(clk_c), 
            .Q(dec_new_block[0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w3_reg__i1.GSR = "ENABLED";
    LUT4 n2757_bdd_4_lut (.A(n2752[27]), .B(n9418), .C(n30146), .D(n25333), 
         .Z(tmp_sboxw[27])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n2757_bdd_4_lut.init = 16'h00ca;
    LUT4 i1_2_lut_3_lut_4_lut (.A(dec_new_block[84]), .B(round_key[84]), 
         .C(n33704), .D(block_new_127__N_1901[69]), .Z(n5)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_451_4_lut (.A(dec_new_block[110]), .B(round_key[110]), 
         .C(dec_new_block[127]), .D(round_key[127]), .Z(n33755)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_rep_451_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_450_4_lut (.A(dec_new_block[109]), .B(round_key[109]), 
         .C(dec_new_block[126]), .D(round_key[126]), .Z(n33754)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_rep_450_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_449_4_lut (.A(dec_new_block[79]), .B(round_key[79]), 
         .C(dec_new_block[95]), .D(round_key[95]), .Z(n33753)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_rep_449_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_448_4_lut (.A(dec_new_block[73]), .B(round_key[73]), 
         .C(dec_new_block[81]), .D(round_key[81]), .Z(n33752)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_448_4_lut.init = 16'h6996;
    FD1P3AX round_ctr_reg_i0_i0 (.D(round_ctr_new[0]), .SP(round_ctr_we), 
            .CK(clk_c), .Q(dec_round_nr[0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam round_ctr_reg_i0_i0.GSR = "ENABLED";
    LUT4 i2_2_lut_3_lut_4_lut (.A(block_new_127__N_1901[67]), .B(n29254), 
         .C(n29172), .D(n29483), .Z(n6)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i2_2_lut_3_lut_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_447_4_lut (.A(dec_new_block[62]), .B(round_key[62]), 
         .C(dec_new_block[54]), .D(round_key[54]), .Z(n33751)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_rep_447_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_446_4_lut (.A(dec_new_block[0]), .B(round_key[0]), 
         .C(dec_new_block[16]), .D(round_key[16]), .Z(n33750)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_rep_446_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_445_4_lut (.A(dec_new_block[31]), .B(round_key[31]), 
         .C(dec_new_block[15]), .D(round_key[15]), .Z(n33749)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_rep_445_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_444_4_lut (.A(dec_new_block[62]), .B(round_key[62]), 
         .C(dec_new_block[41]), .D(round_key[41]), .Z(n33748)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_444_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_220_3_lut (.A(dec_new_block[99]), .B(round_key[99]), 
         .C(n28961), .Z(n33524)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_rep_220_3_lut.init = 16'h9696;
    LUT4 i1_2_lut_rep_202_3_lut (.A(dec_new_block[39]), .B(round_key[39]), 
         .C(n28926), .Z(n33506)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_rep_202_3_lut.init = 16'h9696;
    LUT4 i1_2_lut_4_lut (.A(dec_new_block[117]), .B(round_key[117]), .C(dec_new_block[119]), 
         .D(round_key[119]), .Z(n12084)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_219_3_lut (.A(dec_new_block[3]), .B(round_key[3]), 
         .C(n29447), .Z(n33523)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_rep_219_3_lut.init = 16'h9696;
    LUT4 i1_2_lut_rep_203_3_lut_4_lut (.A(dec_new_block[67]), .B(round_key[67]), 
         .C(n29254), .D(n29483), .Z(n33507)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_rep_203_3_lut_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_218_3_lut (.A(dec_new_block[67]), .B(round_key[67]), 
         .C(n29254), .Z(n33522)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_rep_218_3_lut.init = 16'h9696;
    FD1P3AX block_w1_reg__i1 (.D(n3899[64]), .SP(block_w1_we), .CK(clk_c), 
            .Q(dec_new_block[64])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w1_reg__i1.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i1 (.D(n3899[96]), .SP(block_w0_we), .CK(clk_c), 
            .Q(dec_new_block[96])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w0_reg__i1.GSR = "ENABLED";
    LUT4 n2758_bdd_4_lut (.A(n2752[26]), .B(n9416), .C(n30146), .D(n25333), 
         .Z(tmp_sboxw[26])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n2758_bdd_4_lut.init = 16'h00ca;
    LUT4 i2_4_lut (.A(n6347[3]), .B(n4_c), .C(encdec_reg), .D(\aes_core_ctrl_new_1__N_858[1] ), 
         .Z(n28773)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B)) */ ;
    defparam i2_4_lut.init = 16'hceee;
    LUT4 i1_4_lut (.A(\enc_round_nr[3] ), .B(block_w3_we_N_1490), .C(n4), 
         .D(n6347[1]), .Z(n4_c)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A !(B+!(D))) */ ;
    defparam i1_4_lut.init = 16'hb3a0;
    LUT4 new_block_127__I_0_i125_2_lut (.A(dec_new_block[124]), .B(round_key[124]), 
         .Z(block_new_127__N_1901[124])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i125_2_lut.init = 16'h6666;
    LUT4 i2_3_lut_rep_204_4_lut (.A(block_new_127__N_1901[3]), .B(n29447), 
         .C(n33829), .D(n6228[3]), .Z(n33508)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i2_3_lut_rep_204_4_lut.init = 16'h6996;
    LUT4 i3_3_lut_4_lut (.A(n33673), .B(n33686), .C(block_new_127__N_1901[8]), 
         .D(n33825), .Z(n8)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i3_3_lut_4_lut.init = 16'h6996;
    LUT4 i1_4_lut_adj_59 (.A(dec_round_nr_c[1]), .B(n33858), .C(n149), 
         .D(dec_round_nr[0]), .Z(round_ctr_new_c[1])) /* synthesis lut_function=(A (B+(C (D)))+!A (B+!((D)+!C))) */ ;
    defparam i1_4_lut_adj_59.init = 16'hecdc;
    LUT4 i27545_3_lut_4_lut (.A(block_new_127__N_1645[39]), .B(update_type[0]), 
         .C(n33844), .D(n13131), .Z(n4540[71])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27545_3_lut_4_lut.init = 16'hf808;
    LUT4 i27543_3_lut_4_lut (.A(block_new_127__N_1645_c[38]), .B(update_type[0]), 
         .C(n33844), .D(n13130), .Z(n4540[70])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27543_3_lut_4_lut.init = 16'hf808;
    LUT4 i27693_3_lut_4_lut (.A(\block_new_127__N_1645[37] ), .B(update_type[0]), 
         .C(n33844), .D(n13129), .Z(n4540[69])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27693_3_lut_4_lut.init = 16'hf808;
    LUT4 i27615_3_lut_4_lut (.A(\block_new_127__N_1645[36] ), .B(update_type[0]), 
         .C(n33844), .D(n13128), .Z(n4540[68])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27615_3_lut_4_lut.init = 16'hf808;
    LUT4 i27613_3_lut_4_lut (.A(block_new_127__N_1645_c[35]), .B(update_type[0]), 
         .C(n33844), .D(n13127), .Z(n4540[67])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27613_3_lut_4_lut.init = 16'hf808;
    LUT4 i27611_3_lut_4_lut (.A(\block_new_127__N_1645[34] ), .B(update_type[0]), 
         .C(n33844), .D(n13126), .Z(n4540[66])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27611_3_lut_4_lut.init = 16'hf808;
    LUT4 i27241_3_lut_4_lut (.A(\block_new_127__N_1645[33] ), .B(update_type[0]), 
         .C(n33844), .D(n13125), .Z(n4540[65])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27241_3_lut_4_lut.init = 16'hf808;
    LUT4 i27691_3_lut_4_lut (.A(block_new_127__N_1645_c[32]), .B(update_type[0]), 
         .C(n33844), .D(n13124), .Z(n4540[64])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27691_3_lut_4_lut.init = 16'hf808;
    LUT4 i27541_3_lut_4_lut (.A(block_new_127__N_1645_c[63]), .B(update_type[0]), 
         .C(n33844), .D(n13123), .Z(n4540[63])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27541_3_lut_4_lut.init = 16'hf808;
    LUT4 i3_2_lut_4_lut (.A(n33774), .B(block_new_127__N_1901[10]), .C(block_new_127__N_1901[26]), 
         .D(n33749), .Z(n9)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i3_2_lut_4_lut.init = 16'h6996;
    LUT4 i27539_3_lut_4_lut (.A(\block_new_127__N_1645[62] ), .B(update_type[0]), 
         .C(n33844), .D(n13122), .Z(n4540[62])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27539_3_lut_4_lut.init = 16'hf808;
    LUT4 i27689_3_lut_4_lut (.A(\block_new_127__N_1645[61] ), .B(update_type[0]), 
         .C(n33844), .D(n13121), .Z(n4540[61])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27689_3_lut_4_lut.init = 16'hf808;
    LUT4 i1_2_lut_4_lut_adj_60 (.A(n33679), .B(block_new_127__N_1901[127]), 
         .C(n33766), .D(n33768), .Z(n4_adj_7671)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_4_lut_adj_60.init = 16'h6996;
    LUT4 i27609_3_lut_4_lut (.A(\block_new_127__N_1645[60] ), .B(update_type[0]), 
         .C(n33844), .D(n13120), .Z(n4540[60])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27609_3_lut_4_lut.init = 16'hf808;
    LUT4 n2769_bdd_4_lut (.A(n2752[15]), .B(n9394), .C(n30146), .D(n25333), 
         .Z(tmp_sboxw[15])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n2769_bdd_4_lut.init = 16'h00ca;
    LUT4 i1_2_lut_4_lut_adj_61 (.A(n33675), .B(block_new_127__N_1901[36]), 
         .C(n4770[4]), .D(block_new_127__N_1901[44]), .Z(n4_adj_7672)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_4_lut_adj_61.init = 16'h6996;
    LUT4 i27741_3_lut_4_lut (.A(\block_new_127__N_1645[59] ), .B(update_type[0]), 
         .C(n33844), .D(n13119), .Z(n4540[59])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27741_3_lut_4_lut.init = 16'hf808;
    LUT4 i27239_3_lut_4_lut (.A(block_new_127__N_1645_c[58]), .B(update_type[0]), 
         .C(n33844), .D(n13118), .Z(n4540[58])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27239_3_lut_4_lut.init = 16'hf808;
    LUT4 n2770_bdd_4_lut (.A(n2752[14]), .B(n9392), .C(n30146), .D(n25333), 
         .Z(tmp_sboxw[14])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n2770_bdd_4_lut.init = 16'h00ca;
    LUT4 i3_2_lut_4_lut_adj_62 (.A(n33675), .B(block_new_127__N_1901[36]), 
         .C(n4770[4]), .D(n33751), .Z(n9_adj_7673)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i3_2_lut_4_lut_adj_62.init = 16'h6996;
    LUT4 i27537_3_lut_4_lut (.A(\block_new_127__N_1645[57] ), .B(update_type[0]), 
         .C(n33844), .D(n13117), .Z(n4540[57])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27537_3_lut_4_lut.init = 16'hf808;
    LUT4 i27535_3_lut_4_lut (.A(block_new_127__N_1645_c[56]), .B(update_type[0]), 
         .C(n33844), .D(n13116), .Z(n4540[56])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27535_3_lut_4_lut.init = 16'hf808;
    LUT4 n2759_bdd_4_lut (.A(n2752[25]), .B(n9414), .C(n30146), .D(n25333), 
         .Z(tmp_sboxw[25])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n2759_bdd_4_lut.init = 16'h00ca;
    LUT4 n2771_bdd_4_lut (.A(n2752[13]), .B(n9390), .C(n30146), .D(n25333), 
         .Z(tmp_sboxw[13])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n2771_bdd_4_lut.init = 16'h00ca;
    LUT4 i2_2_lut_4_lut (.A(n33675), .B(block_new_127__N_1901[36]), .C(n4770[4]), 
         .D(block_new_127__N_1901[38]), .Z(n7)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i2_2_lut_4_lut.init = 16'h6996;
    LUT4 i27237_3_lut_4_lut (.A(\block_new_127__N_1645[87] ), .B(update_type[0]), 
         .C(n33844), .D(n13115), .Z(n4540[55])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27237_3_lut_4_lut.init = 16'hf808;
    LUT4 i3_3_lut_4_lut_adj_63 (.A(block_new_127__N_1901[99]), .B(n28961), 
         .C(block_new_127__N_1901[123]), .D(n29441), .Z(n8_adj_7674)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i3_3_lut_4_lut_adj_63.init = 16'h6996;
    LUT4 i2_3_lut_rep_205_4_lut (.A(block_new_127__N_1901[99]), .B(n28961), 
         .C(n873[3]), .D(n648[3]), .Z(n33509)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i2_3_lut_rep_205_4_lut.init = 16'h6996;
    LUT4 n2772_bdd_4_lut (.A(n2752[12]), .B(n9388), .C(n30146), .D(n25333), 
         .Z(tmp_sboxw[12])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n2772_bdd_4_lut.init = 16'h00ca;
    LUT4 i3_2_lut_3_lut_4_lut (.A(block_new_127__N_1901[88]), .B(n33796), 
         .C(n33752), .D(n33803), .Z(n9_adj_7675)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i3_2_lut_3_lut_4_lut.init = 16'h6996;
    LUT4 i27533_3_lut_4_lut (.A(\block_new_127__N_1645[86] ), .B(update_type[0]), 
         .C(n33844), .D(n13114), .Z(n4540[54])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27533_3_lut_4_lut.init = 16'hf808;
    LUT4 n2773_bdd_4_lut (.A(n2752[11]), .B(n9386), .C(n30146), .D(n25333), 
         .Z(tmp_sboxw[11])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n2773_bdd_4_lut.init = 16'h00ca;
    LUT4 i27687_3_lut_4_lut (.A(\block_new_127__N_1645[85] ), .B(update_type[0]), 
         .C(n33844), .D(n13113), .Z(n4540[53])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27687_3_lut_4_lut.init = 16'hf808;
    LUT4 i27685_3_lut_4_lut (.A(\block_new_127__N_1645[84] ), .B(update_type[0]), 
         .C(n33844), .D(n13112), .Z(n4540[52])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27685_3_lut_4_lut.init = 16'hf808;
    LUT4 n2774_bdd_4_lut (.A(n2752[10]), .B(n9384), .C(n30146), .D(n25333), 
         .Z(tmp_sboxw[10])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n2774_bdd_4_lut.init = 16'h00ca;
    LUT4 n2775_bdd_4_lut (.A(n2752[9]), .B(n9382), .C(n30146), .D(n25333), 
         .Z(tmp_sboxw[9])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n2775_bdd_4_lut.init = 16'h00ca;
    LUT4 i3_3_lut_4_lut_adj_64 (.A(block_new_127__N_1901[39]), .B(n28926), 
         .C(block_new_127__N_1901[63]), .D(block_new_127__N_1901[32]), .Z(n8_adj_7676)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i3_3_lut_4_lut_adj_64.init = 16'h6996;
    LUT4 n2776_bdd_4_lut (.A(n2752[8]), .B(n9380), .C(n30146), .D(n25333), 
         .Z(tmp_sboxw[8])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n2776_bdd_4_lut.init = 16'h00ca;
    LUT4 i2_2_lut_4_lut_adj_65 (.A(block_new_127__N_1901[105]), .B(block_new_127__N_1901[110]), 
         .C(n33678), .D(n33688), .Z(n7_adj_7677)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i2_2_lut_4_lut_adj_65.init = 16'h6996;
    LUT4 i2_2_lut_4_lut_adj_66 (.A(n33804), .B(block_new_127__N_1901[87]), 
         .C(block_new_127__N_1901[64]), .D(n33681), .Z(n7_adj_7678)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i2_2_lut_4_lut_adj_66.init = 16'h6996;
    LUT4 i2_2_lut_4_lut_adj_67 (.A(n33692), .B(n33702), .C(n33796), .D(block_new_127__N_1901[85]), 
         .Z(n6_adj_7679)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i2_2_lut_4_lut_adj_67.init = 16'h6996;
    LUT4 n2760_bdd_4_lut (.A(n2752[24]), .B(n9412), .C(n30146), .D(n25333), 
         .Z(tmp_sboxw[24])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n2760_bdd_4_lut.init = 16'h00ca;
    LUT4 i27789_3_lut_4_lut (.A(\block_new_127__N_1645[83] ), .B(update_type[0]), 
         .C(n33844), .D(n13111), .Z(n4540[51])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27789_3_lut_4_lut.init = 16'hf808;
    LUT4 i27531_3_lut_4_lut (.A(\block_new_127__N_1645[82] ), .B(update_type[0]), 
         .C(n33844), .D(n13110), .Z(n4540[50])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27531_3_lut_4_lut.init = 16'hf808;
    LUT4 i1_2_lut_4_lut_adj_68 (.A(n33804), .B(block_new_127__N_1901[87]), 
         .C(block_new_127__N_1901[64]), .D(n33820), .Z(n4_adj_7680)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_4_lut_adj_68.init = 16'h6996;
    LUT4 n2777_bdd_4_lut (.A(n2752[7]), .B(n9378), .C(n30146), .D(n25333), 
         .Z(tmp_sboxw[7])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n2777_bdd_4_lut.init = 16'h00ca;
    LUT4 i27739_3_lut_4_lut (.A(\block_new_127__N_1645[81] ), .B(update_type[0]), 
         .C(n33844), .D(n13109), .Z(n4540[49])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27739_3_lut_4_lut.init = 16'hf808;
    LUT4 i1_2_lut_4_lut_adj_69 (.A(n33692), .B(n33702), .C(n33796), .D(block_new_127__N_1901[77]), 
         .Z(n5_adj_7681)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_4_lut_adj_69.init = 16'h6996;
    LUT4 i27235_3_lut_4_lut (.A(block_new_127__N_1645_c[80]), .B(update_type[0]), 
         .C(n33844), .D(n13108), .Z(n4540[48])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27235_3_lut_4_lut.init = 16'hf808;
    LUT4 i27607_3_lut_4_lut (.A(block_new_127__N_1645_c[111]), .B(update_type[0]), 
         .C(n33844), .D(n13107), .Z(n4540[47])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27607_3_lut_4_lut.init = 16'hf808;
    LUT4 i27529_3_lut_4_lut (.A(block_new_127__N_1645_c[110]), .B(update_type[0]), 
         .C(n33844), .D(n13106), .Z(n4540[46])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27529_3_lut_4_lut.init = 16'hf808;
    LUT4 n2778_bdd_4_lut (.A(n2752[6]), .B(n9376), .C(n30146), .D(n25333), 
         .Z(tmp_sboxw[6])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n2778_bdd_4_lut.init = 16'h00ca;
    LUT4 i27683_3_lut_4_lut (.A(block_new_127__N_1645_c[109]), .B(update_type[0]), 
         .C(n33844), .D(n13105), .Z(n4540[45])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27683_3_lut_4_lut.init = 16'hf808;
    LUT4 i3_3_lut_4_lut_adj_70 (.A(block_new_127__N_1901[93]), .B(n33683), 
         .C(n33703), .D(n29381), .Z(n8_adj_7682)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i3_3_lut_4_lut_adj_70.init = 16'h6996;
    LUT4 i2_2_lut_3_lut_4_lut_adj_71 (.A(n33804), .B(n33785), .C(n33753), 
         .D(n33794), .Z(n6_adj_7683)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i2_2_lut_3_lut_4_lut_adj_71.init = 16'h6996;
    LUT4 n2779_bdd_4_lut (.A(n2752[5]), .B(n9374), .C(n30146), .D(n25333), 
         .Z(tmp_sboxw[5])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n2779_bdd_4_lut.init = 16'h00ca;
    LUT4 i27681_3_lut_4_lut (.A(\block_new_127__N_1645[108] ), .B(update_type[0]), 
         .C(n33844), .D(n13104), .Z(n4540[44])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27681_3_lut_4_lut.init = 16'hf808;
    LUT4 n2780_bdd_4_lut (.A(n2752[4]), .B(n9372), .C(n30146), .D(n25333), 
         .Z(tmp_sboxw[4])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n2780_bdd_4_lut.init = 16'h00ca;
    LUT4 i27737_3_lut_4_lut (.A(\block_new_127__N_1645[107] ), .B(update_type[0]), 
         .C(n33844), .D(n13103), .Z(n4540[43])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27737_3_lut_4_lut.init = 16'hf808;
    LUT4 i27605_3_lut_4_lut (.A(block_new_127__N_1645_c[106]), .B(update_type[0]), 
         .C(n33844), .D(n13102), .Z(n4540[42])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27605_3_lut_4_lut.init = 16'hf808;
    LUT4 n2781_bdd_4_lut (.A(n2752[3]), .B(n9370), .C(n30146), .D(n25333), 
         .Z(tmp_sboxw[3])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n2781_bdd_4_lut.init = 16'h00ca;
    LUT4 i3_3_lut_4_lut_adj_72 (.A(n4770[4]), .B(n33699), .C(n33706), 
         .D(n33684), .Z(n8_adj_7684)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i3_3_lut_4_lut_adj_72.init = 16'h6996;
    LUT4 i27603_3_lut_4_lut (.A(\block_new_127__N_1645[105] ), .B(update_type[0]), 
         .C(n33844), .D(n13101), .Z(n4540[41])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27603_3_lut_4_lut.init = 16'hf808;
    LUT4 i27527_3_lut_4_lut (.A(block_new_127__N_1645_c[104]), .B(update_type[0]), 
         .C(n33844), .D(n13100), .Z(n4540[40])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27527_3_lut_4_lut.init = 16'hf808;
    LUT4 i27525_3_lut_4_lut (.A(\block_new_127__N_1645[7] ), .B(update_type[0]), 
         .C(n33844), .D(n13099), .Z(n4540[39])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27525_3_lut_4_lut.init = 16'hf808;
    LUT4 i27601_3_lut_4_lut (.A(block_new_127__N_1645_c[6]), .B(update_type[0]), 
         .C(n33844), .D(n13098), .Z(n4540[38])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27601_3_lut_4_lut.init = 16'hf808;
    LUT4 n2782_bdd_4_lut (.A(n2752[2]), .B(n9368), .C(n30146), .D(n25333), 
         .Z(tmp_sboxw[2])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n2782_bdd_4_lut.init = 16'h00ca;
    LUT4 i27599_3_lut_4_lut (.A(\block_new_127__N_1645[5] ), .B(update_type[0]), 
         .C(n33844), .D(n13097), .Z(n4540[37])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27599_3_lut_4_lut.init = 16'hf808;
    LUT4 i2_2_lut_3_lut_4_lut_adj_73 (.A(block_new_127__N_1901[53]), .B(n33801), 
         .C(n33772), .D(block_new_127__N_1901[48]), .Z(n6_adj_7685)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i2_2_lut_3_lut_4_lut_adj_73.init = 16'h6996;
    LUT4 i27679_3_lut_4_lut (.A(\block_new_127__N_1645[4] ), .B(update_type[0]), 
         .C(n33844), .D(n13096), .Z(n4540[36])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27679_3_lut_4_lut.init = 16'hf808;
    LUT4 i27677_3_lut_4_lut (.A(\block_new_127__N_1645[3] ), .B(update_type[0]), 
         .C(n33844), .D(n13095), .Z(n4540[35])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27677_3_lut_4_lut.init = 16'hf808;
    LUT4 i3_3_lut_4_lut_adj_74 (.A(block_new_127__N_1901[53]), .B(n33801), 
         .C(block_new_127__N_1901[45]), .D(n33707), .Z(n8_adj_7686)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i3_3_lut_4_lut_adj_74.init = 16'h6996;
    LUT4 i27523_3_lut_4_lut (.A(\block_new_127__N_1645[2] ), .B(update_type[0]), 
         .C(n33844), .D(n13094), .Z(n4540[34])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27523_3_lut_4_lut.init = 16'hf808;
    LUT4 i9396_3_lut (.A(dec_round_nr_c[1]), .B(\enc_round_nr[1] ), .C(encdec_reg), 
         .Z(\muxed_round_nr[1] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(96[7:17])
    defparam i9396_3_lut.init = 16'hcaca;
    LUT4 i3_3_lut_4_lut_adj_75 (.A(block_new_127__N_1901[105]), .B(n33689), 
         .C(block_new_127__N_1901[97]), .D(block_new_127__N_1901[112]), 
         .Z(n8_adj_7687)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i3_3_lut_4_lut_adj_75.init = 16'h6996;
    LUT4 i3_3_lut_4_lut_adj_76 (.A(n33836), .B(n29160), .C(n33838), .D(block_new_127__N_1901[101]), 
         .Z(n8_adj_7688)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i3_3_lut_4_lut_adj_76.init = 16'h6996;
    LUT4 i27675_3_lut_4_lut (.A(\block_new_127__N_1645[1] ), .B(update_type[0]), 
         .C(n33844), .D(n13093), .Z(n4540[33])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27675_3_lut_4_lut.init = 16'hf808;
    LUT4 i27521_3_lut_4_lut (.A(block_new_127__N_1645_c[0]), .B(update_type[0]), 
         .C(n33844), .D(n13092), .Z(n4540[32])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27521_3_lut_4_lut.init = 16'hf808;
    LUT4 n2783_bdd_4_lut (.A(n2752[1]), .B(n9366), .C(n30146), .D(n25333), 
         .Z(tmp_sboxw[1])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n2783_bdd_4_lut.init = 16'h00ca;
    LUT4 n2784_bdd_4_lut (.A(n2752[0]), .B(n8522), .C(n30146), .D(n25333), 
         .Z(tmp_sboxw[0])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n2784_bdd_4_lut.init = 16'h00ca;
    LUT4 i2_2_lut_4_lut_adj_77 (.A(n33763), .B(n33800), .C(n33685), .D(block_new_127__N_1901[63]), 
         .Z(n6_adj_7689)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i2_2_lut_4_lut_adj_77.init = 16'h6996;
    LUT4 i4_3_lut_4_lut (.A(block_new_127__N_1901[62]), .B(n33786), .C(block_new_127__N_1901[41]), 
         .D(block_new_127__N_1901[58]), .Z(n11)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i4_3_lut_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_3_lut (.A(block_new_127__N_1901[62]), .B(block_new_127__N_1901[41]), 
         .C(n28987), .Z(n4_adj_7690)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_3_lut.init = 16'h9696;
    LUT4 i2_2_lut_3_lut_4_lut_adj_78 (.A(n33754), .B(n33755), .C(n33689), 
         .D(block_new_127__N_1901[105]), .Z(n6_adj_7691)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i2_2_lut_3_lut_4_lut_adj_78.init = 16'h6996;
    LUT4 i1_2_lut_3_lut_4_lut_adj_79 (.A(block_new_127__N_1901[62]), .B(block_new_127__N_1901[41]), 
         .C(n33813), .D(block_new_127__N_1901[57]), .Z(n5_adj_7692)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_3_lut_4_lut_adj_79.init = 16'h6996;
    LUT4 i27597_3_lut_4_lut (.A(block_new_127__N_1645_c[31]), .B(update_type[0]), 
         .C(n33844), .D(n13091), .Z(n4540[31])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27597_3_lut_4_lut.init = 16'hf808;
    LUT4 i2_2_lut_3_lut_4_lut_adj_80 (.A(n33791), .B(n33756), .C(n33755), 
         .D(n33754), .Z(n6_adj_7693)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i2_2_lut_3_lut_4_lut_adj_80.init = 16'h6996;
    LUT4 i27595_3_lut_4_lut (.A(\block_new_127__N_1645[30] ), .B(update_type[0]), 
         .C(n33844), .D(n13090), .Z(n4540[30])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27595_3_lut_4_lut.init = 16'hf808;
    LUT4 n2761_bdd_4_lut (.A(n2752[23]), .B(n9410), .C(n30146), .D(n25333), 
         .Z(tmp_sboxw[23])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n2761_bdd_4_lut.init = 16'h00ca;
    LUT4 i3_3_lut_4_lut_adj_81 (.A(n33791), .B(n33756), .C(block_new_127__N_1901[111]), 
         .D(block_new_127__N_1901[120]), .Z(n8_adj_7694)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i3_3_lut_4_lut_adj_81.init = 16'h6996;
    LUT4 mux_626_Mux_1_i2_4_lut (.A(new_sboxw[1]), .B(n5_adj_7695), .C(update_type[0]), 
         .D(n6_adj_7691), .Z(n2)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_1_i2_4_lut.init = 16'h3aca;
    LUT4 mux_626_Mux_13_i2_4_lut (.A(new_sboxw[13]), .B(n5_adj_7696), .C(update_type[0]), 
         .D(n6_adj_7697), .Z(n2_adj_7698)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_13_i2_4_lut.init = 16'h3aca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_82 (.A(block_new_127__N_1901[31]), .B(block_new_127__N_1901[15]), 
         .C(n33774), .D(block_new_127__N_1901[7]), .Z(n4_adj_7699)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_3_lut_4_lut_adj_82.init = 16'h6996;
    LUT4 mux_626_Mux_15_i2_4_lut (.A(new_sboxw[15]), .B(n7_adj_7700), .C(update_type[0]), 
         .D(n8_adj_7701), .Z(n2_adj_7702)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_15_i2_4_lut.init = 16'h3aca;
    LUT4 mux_626_Mux_17_i2_4_lut (.A(new_sboxw[17]), .B(n5_adj_7692), .C(update_type[0]), 
         .D(n6_adj_7703), .Z(n2_adj_7704)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_17_i2_4_lut.init = 16'h3aca;
    LUT4 mux_626_Mux_18_i2_4_lut (.A(new_sboxw[18]), .B(n29390), .C(update_type[0]), 
         .D(n4_adj_7690), .Z(n2_adj_7705)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_18_i2_4_lut.init = 16'h3aca;
    LUT4 mux_626_Mux_22_i2_4_lut (.A(new_sboxw[22]), .B(n7), .C(update_type[0]), 
         .D(n8_adj_7686), .Z(n2_adj_7706)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_22_i2_4_lut.init = 16'h3aca;
    LUT4 mux_626_Mux_25_i2_4_lut (.A(new_sboxw[25]), .B(n9_adj_7707), .C(update_type[0]), 
         .D(n10), .Z(n2_adj_7708)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_25_i2_4_lut.init = 16'h3aca;
    LUT4 i2_3_lut_rep_214_4_lut (.A(n33688), .B(block_new_127__N_1901[106]), 
         .C(block_new_127__N_1901[114]), .D(block_new_127__N_1901[121]), 
         .Z(n33518)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i2_3_lut_rep_214_4_lut.init = 16'h6996;
    LUT4 mux_626_Mux_32_i2_4_lut (.A(new_sboxw[0]), .B(n7_adj_7709), .C(update_type[0]), 
         .D(n8), .Z(n2_adj_7710)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_32_i2_4_lut.init = 16'h3aca;
    LUT4 mux_626_Mux_34_i2_4_lut (.A(new_sboxw[2]), .B(n9), .C(update_type[0]), 
         .D(n10_adj_7711), .Z(n2_adj_7712)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_34_i2_4_lut.init = 16'h3aca;
    LUT4 mux_626_Mux_39_i2_4_lut (.A(new_sboxw[7]), .B(n5_adj_7713), .C(update_type[0]), 
         .D(n6_adj_7714), .Z(n2_adj_7715)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_39_i2_4_lut.init = 16'h3aca;
    LUT4 mux_626_Mux_40_i2_4_lut (.A(new_sboxw[8]), .B(n7_adj_7716), .C(update_type[0]), 
         .D(n8_adj_7694), .Z(n2_adj_7717)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_40_i2_4_lut.init = 16'h3aca;
    LUT4 i3_3_lut_4_lut_adj_83 (.A(block_new_127__N_1901[117]), .B(n33690), 
         .C(block_new_127__N_1901[124]), .D(n33589), .Z(n8_adj_7718)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i3_3_lut_4_lut_adj_83.init = 16'h6996;
    LUT4 mux_626_Mux_46_i2_4_lut (.A(new_sboxw[14]), .B(n5_adj_7719), .C(update_type[0]), 
         .D(n6_adj_7720), .Z(n2_adj_7721)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_46_i2_4_lut.init = 16'h3aca;
    LUT4 mux_626_Mux_50_i2_4_lut (.A(new_sboxw[18]), .B(n29396), .C(update_type[0]), 
         .D(n4_adj_7722), .Z(n2_adj_7723)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_50_i2_4_lut.init = 16'h3aca;
    LUT4 mux_626_Mux_54_i2_4_lut (.A(new_sboxw[22]), .B(n7_adj_7724), .C(update_type[0]), 
         .D(n8_adj_7725), .Z(n2_adj_7726)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_54_i2_4_lut.init = 16'h3aca;
    LUT4 mux_626_Mux_56_i2_4_lut (.A(new_sboxw[24]), .B(n7_adj_7727), .C(update_type[0]), 
         .D(n8_adj_7728), .Z(n2_adj_7729)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_56_i2_4_lut.init = 16'h3aca;
    LUT4 i2_2_lut_3_lut_4_lut_adj_84 (.A(block_new_127__N_1901[0]), .B(block_new_127__N_1901[16]), 
         .C(n33781), .D(n33757), .Z(n7_adj_7730)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i2_2_lut_3_lut_4_lut_adj_84.init = 16'h6996;
    LUT4 i27673_3_lut_4_lut (.A(block_new_127__N_1645_c[29]), .B(update_type[0]), 
         .C(n33844), .D(n13089), .Z(n4540[29])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27673_3_lut_4_lut.init = 16'hf808;
    LUT4 i27671_3_lut_4_lut (.A(\block_new_127__N_1645[28] ), .B(update_type[0]), 
         .C(n33844), .D(n13088), .Z(n4540[28])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27671_3_lut_4_lut.init = 16'hf808;
    LUT4 i3_3_lut_4_lut_adj_85 (.A(block_new_127__N_1901[117]), .B(n33690), 
         .C(n33710), .D(n33839), .Z(n8_adj_7731)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i3_3_lut_4_lut_adj_85.init = 16'h6996;
    LUT4 mux_626_Mux_57_i2_4_lut (.A(new_sboxw[25]), .B(n7_adj_7732), .C(update_type[0]), 
         .D(n8_adj_7733), .Z(n2_adj_7734)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_57_i2_4_lut.init = 16'h3aca;
    LUT4 mux_626_Mux_62_i2_4_lut (.A(new_sboxw[30]), .B(n9_adj_7735), .C(update_type[0]), 
         .D(n10_adj_7736), .Z(n2_adj_7737)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_62_i2_4_lut.init = 16'h3aca;
    LUT4 i27787_3_lut_4_lut (.A(\block_new_127__N_1645[27] ), .B(update_type[0]), 
         .C(n33844), .D(n13087), .Z(n4540[27])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27787_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_626_Mux_63_i2_4_lut (.A(new_sboxw[31]), .B(n33582), .C(update_type[0]), 
         .D(n4_adj_7738), .Z(n2_adj_7739)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_63_i2_4_lut.init = 16'h3aca;
    LUT4 i27669_3_lut_4_lut (.A(block_new_127__N_1645_c[26]), .B(update_type[0]), 
         .C(n33844), .D(n13086), .Z(n4540[26])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27669_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_626_Mux_70_i2_4_lut (.A(new_sboxw[6]), .B(n9_adj_7673), .C(update_type[0]), 
         .D(n10_adj_7740), .Z(n2_adj_7741)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_70_i2_4_lut.init = 16'h3aca;
    LUT4 i27519_3_lut_4_lut (.A(\block_new_127__N_1645[25] ), .B(update_type[0]), 
         .C(n33844), .D(n13085), .Z(n4540[25])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27519_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_626_Mux_71_i2_4_lut (.A(new_sboxw[7]), .B(n5_adj_7742), .C(update_type[0]), 
         .D(n6_adj_7743), .Z(n2_adj_7744)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_71_i2_4_lut.init = 16'h3aca;
    LUT4 mux_626_Mux_73_i2_4_lut (.A(new_sboxw[9]), .B(n9_adj_7745), .C(update_type[0]), 
         .D(n10_adj_7746), .Z(n2_adj_7747)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_73_i2_4_lut.init = 16'h3aca;
    LUT4 mux_626_Mux_79_i2_4_lut (.A(new_sboxw[15]), .B(n33580), .C(update_type[0]), 
         .D(n4_adj_7748), .Z(n2_adj_7749)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_79_i2_4_lut.init = 16'h3aca;
    LUT4 i27667_3_lut_4_lut (.A(block_new_127__N_1645_c[24]), .B(update_type[0]), 
         .C(n33844), .D(n13084), .Z(n4540[24])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27667_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_626_Mux_80_i2_4_lut (.A(new_sboxw[16]), .B(n29375), .C(update_type[0]), 
         .D(n4_adj_7750), .Z(n2_adj_7751)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_80_i2_4_lut.init = 16'h3aca;
    LUT4 new_block_127__I_0_i124_2_lut (.A(dec_new_block[123]), .B(round_key[123]), 
         .Z(block_new_127__N_1901[123])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i124_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i123_2_lut (.A(\block_reg[0] [26]), .B(round_key[122]), 
         .Z(block_new_127__N_1645_c[122])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i123_2_lut.init = 16'h6666;
    LUT4 i1_2_lut_3_lut_adj_86 (.A(block_new_127__N_1901[62]), .B(block_new_127__N_1901[54]), 
         .C(n28987), .Z(n5_adj_7752)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_3_lut_adj_86.init = 16'h9696;
    LUT4 i3081_3_lut (.A(dec_new_block[32]), .B(dec_new_block[0]), .C(n6362[3]), 
         .Z(n8522)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam i3081_3_lut.init = 16'hcaca;
    LUT4 mux_626_Mux_82_i2_4_lut (.A(new_sboxw[18]), .B(n7_adj_7753), .C(update_type[0]), 
         .D(n8_adj_7754), .Z(n2_adj_7755)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_82_i2_4_lut.init = 16'h3aca;
    LUT4 mux_224_i1_3_lut (.A(dec_new_block[96]), .B(dec_new_block[64]), 
         .C(n6362[1]), .Z(n2752[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam mux_224_i1_3_lut.init = 16'hcaca;
    LUT4 i27233_3_lut_4_lut (.A(block_new_127__N_1645_c[55]), .B(update_type[0]), 
         .C(n33844), .D(n13083), .Z(n4540[23])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27233_3_lut_4_lut.init = 16'hf808;
    LUT4 i27517_3_lut_4_lut (.A(block_new_127__N_1645_c[54]), .B(update_type[0]), 
         .C(n33844), .D(n13082), .Z(n4540[22])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27517_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_626_Mux_86_i2_4_lut (.A(new_sboxw[22]), .B(n7_adj_7756), .C(update_type[0]), 
         .D(n8_adj_7731), .Z(n2_adj_7757)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_86_i2_4_lut.init = 16'h3aca;
    LUT4 i3757_3_lut (.A(dec_new_block[33]), .B(dec_new_block[1]), .C(n6362[3]), 
         .Z(n9366)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam i3757_3_lut.init = 16'hcaca;
    LUT4 mux_224_i2_3_lut (.A(dec_new_block[97]), .B(dec_new_block[65]), 
         .C(n6362[1]), .Z(n2752[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam mux_224_i2_3_lut.init = 16'hcaca;
    LUT4 i3759_3_lut (.A(dec_new_block[34]), .B(dec_new_block[2]), .C(n6362[3]), 
         .Z(n9368)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam i3759_3_lut.init = 16'hcaca;
    LUT4 mux_224_i3_3_lut (.A(dec_new_block[98]), .B(dec_new_block[66]), 
         .C(n6362[1]), .Z(n2752[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam mux_224_i3_3_lut.init = 16'hcaca;
    LUT4 i3_3_lut_4_lut_adj_87 (.A(block_new_127__N_1901[31]), .B(block_new_127__N_1901[6]), 
         .C(block_new_127__N_1901[2]), .D(n33668), .Z(n8_adj_7758)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i3_3_lut_4_lut_adj_87.init = 16'h6996;
    LUT4 mux_626_Mux_89_i2_4_lut (.A(new_sboxw[25]), .B(n9_adj_7675), .C(update_type[0]), 
         .D(n10_adj_7759), .Z(n2_adj_7760)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_89_i2_4_lut.init = 16'h3aca;
    LUT4 i3761_3_lut (.A(dec_new_block[35]), .B(dec_new_block[3]), .C(n6362[3]), 
         .Z(n9370)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam i3761_3_lut.init = 16'hcaca;
    LUT4 mux_224_i4_3_lut (.A(dec_new_block[99]), .B(dec_new_block[67]), 
         .C(n6362[1]), .Z(n2752[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam mux_224_i4_3_lut.init = 16'hcaca;
    LUT4 mux_626_Mux_96_i2_4_lut (.A(new_sboxw[0]), .B(n5_adj_7761), .C(update_type[0]), 
         .D(n6_adj_7762), .Z(n2_adj_7763)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_96_i2_4_lut.init = 16'h3aca;
    LUT4 i3763_3_lut (.A(dec_new_block[36]), .B(dec_new_block[4]), .C(n6362[3]), 
         .Z(n9372)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam i3763_3_lut.init = 16'hcaca;
    LUT4 mux_224_i5_3_lut (.A(dec_new_block[100]), .B(dec_new_block[68]), 
         .C(n6362[1]), .Z(n2752[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam mux_224_i5_3_lut.init = 16'hcaca;
    LUT4 i2_2_lut_3_lut_4_lut_adj_88 (.A(block_new_127__N_1901[31]), .B(block_new_127__N_1901[6]), 
         .C(n33677), .D(n12090), .Z(n6_adj_7714)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i2_2_lut_3_lut_4_lut_adj_88.init = 16'h6996;
    LUT4 i3765_3_lut (.A(dec_new_block[37]), .B(dec_new_block[5]), .C(n6362[3]), 
         .Z(n9374)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam i3765_3_lut.init = 16'hcaca;
    LUT4 mux_224_i6_3_lut (.A(dec_new_block[101]), .B(dec_new_block[69]), 
         .C(n6362[1]), .Z(n2752[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam mux_224_i6_3_lut.init = 16'hcaca;
    LUT4 i27593_3_lut_4_lut (.A(block_new_127__N_1645_c[53]), .B(update_type[0]), 
         .C(n33844), .D(n13081), .Z(n4540[21])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27593_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_626_Mux_97_i2_4_lut (.A(new_sboxw[1]), .B(n7_adj_7678), .C(update_type[0]), 
         .D(n8_adj_7764), .Z(n2_adj_7765)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_97_i2_4_lut.init = 16'h3aca;
    LUT4 i3767_3_lut (.A(dec_new_block[38]), .B(dec_new_block[6]), .C(n6362[3]), 
         .Z(n9376)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam i3767_3_lut.init = 16'hcaca;
    LUT4 mux_224_i7_3_lut (.A(dec_new_block[102]), .B(dec_new_block[70]), 
         .C(n6362[1]), .Z(n2752[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam mux_224_i7_3_lut.init = 16'hcaca;
    LUT4 i27591_3_lut_4_lut (.A(block_new_127__N_1645_c[52]), .B(update_type[0]), 
         .C(n33844), .D(n13080), .Z(n4540[20])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27591_3_lut_4_lut.init = 16'hf808;
    LUT4 i27665_3_lut_4_lut (.A(\block_new_127__N_1645[51] ), .B(update_type[0]), 
         .C(n33844), .D(n13079), .Z(n4540[19])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27665_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_626_Mux_98_i2_4_lut (.A(new_sboxw[2]), .B(n29396), .C(update_type[0]), 
         .D(n4_adj_7766), .Z(n2_adj_7767)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_98_i2_4_lut.init = 16'h3aca;
    LUT4 i3769_3_lut (.A(dec_new_block[39]), .B(dec_new_block[7]), .C(n6362[3]), 
         .Z(n9378)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam i3769_3_lut.init = 16'hcaca;
    LUT4 mux_224_i8_3_lut (.A(dec_new_block[103]), .B(dec_new_block[71]), 
         .C(n6362[1]), .Z(n2752[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam mux_224_i8_3_lut.init = 16'hcaca;
    LUT4 i27515_3_lut_4_lut (.A(\block_new_127__N_1645[50] ), .B(update_type[0]), 
         .C(n33844), .D(n13078), .Z(n4540[18])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27515_3_lut_4_lut.init = 16'hf808;
    LUT4 i3771_3_lut (.A(dec_new_block[40]), .B(dec_new_block[8]), .C(n6362[3]), 
         .Z(n9380)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam i3771_3_lut.init = 16'hcaca;
    LUT4 new_block_127__I_0_i109_2_lut (.A(dec_new_block[108]), .B(round_key[108]), 
         .Z(block_new_127__N_1901[108])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i109_2_lut.init = 16'h6666;
    LUT4 i2_2_lut_4_lut_adj_89 (.A(n33523), .B(n6228[3]), .C(n33829), 
         .D(n33713), .Z(n6_adj_7768)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i2_2_lut_4_lut_adj_89.init = 16'h6996;
    LUT4 n2762_bdd_4_lut (.A(n2752[22]), .B(n9408), .C(n30146), .D(n25333), 
         .Z(tmp_sboxw[22])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n2762_bdd_4_lut.init = 16'h00ca;
    LUT4 i3_3_lut_4_lut_adj_90 (.A(block_new_127__N_1901[73]), .B(block_new_127__N_1901[81]), 
         .C(n3564[3]), .D(block_new_127__N_1901[89]), .Z(n8_adj_7764)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i3_3_lut_4_lut_adj_90.init = 16'h6996;
    LUT4 mux_626_Mux_103_i2_4_lut (.A(new_sboxw[7]), .B(n5_adj_7769), .C(update_type[0]), 
         .D(n6_adj_7683), .Z(n2_adj_7770)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_103_i2_4_lut.init = 16'h3aca;
    LUT4 new_block_127__I_0_i102_2_lut (.A(dec_new_block[101]), .B(round_key[101]), 
         .Z(block_new_127__N_1901[101])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i102_2_lut.init = 16'h6666;
    LUT4 mux_626_Mux_104_i2_4_lut (.A(new_sboxw[8]), .B(n5_adj_7771), .C(update_type[0]), 
         .D(n6_adj_7685), .Z(n2_adj_7772)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_104_i2_4_lut.init = 16'h3aca;
    LUT4 mux_224_i9_3_lut (.A(dec_new_block[104]), .B(dec_new_block[72]), 
         .C(n6362[1]), .Z(n2752[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam mux_224_i9_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_adj_91 (.A(block_new_127__N_1901[73]), .B(block_new_127__N_1901[81]), 
         .C(block_new_127__N_1901[66]), .Z(n4_adj_7722)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_3_lut_adj_91.init = 16'h9696;
    LUT4 i3773_3_lut (.A(dec_new_block[41]), .B(dec_new_block[9]), .C(n6362[3]), 
         .Z(n9382)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam i3773_3_lut.init = 16'hcaca;
    LUT4 mux_626_Mux_106_i2_4_lut (.A(new_sboxw[10]), .B(n11), .C(update_type[0]), 
         .D(n12), .Z(n2_adj_7773)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_106_i2_4_lut.init = 16'h3aca;
    LUT4 mux_224_i10_3_lut (.A(dec_new_block[105]), .B(dec_new_block[73]), 
         .C(n6362[1]), .Z(n2752[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam mux_224_i10_3_lut.init = 16'hcaca;
    LUT4 mux_626_Mux_110_i2_4_lut (.A(new_sboxw[14]), .B(n5_adj_7774), .C(update_type[0]), 
         .D(n6_adj_7775), .Z(n2_adj_7776)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_110_i2_4_lut.init = 16'h3aca;
    LUT4 i3775_3_lut (.A(dec_new_block[42]), .B(dec_new_block[10]), .C(n6362[3]), 
         .Z(n9384)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam i3775_3_lut.init = 16'hcaca;
    LUT4 i27513_3_lut_4_lut (.A(\block_new_127__N_1645[49] ), .B(update_type[0]), 
         .C(n33844), .D(n13077), .Z(n4540[17])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27513_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_626_Mux_112_i2_4_lut (.A(new_sboxw[16]), .B(n5_adj_7777), .C(update_type[0]), 
         .D(n6_adj_7778), .Z(n2_adj_7779)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_112_i2_4_lut.init = 16'h3aca;
    LUT4 mux_224_i11_3_lut (.A(dec_new_block[106]), .B(dec_new_block[74]), 
         .C(n6362[1]), .Z(n2752[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam mux_224_i11_3_lut.init = 16'hcaca;
    LUT4 i3777_3_lut (.A(dec_new_block[43]), .B(dec_new_block[11]), .C(n6362[3]), 
         .Z(n9386)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam i3777_3_lut.init = 16'hcaca;
    LUT4 mux_626_Mux_120_i2_4_lut (.A(new_sboxw[24]), .B(n5_adj_7780), .C(update_type[0]), 
         .D(n6_adj_7693), .Z(n2_adj_7781)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_120_i2_4_lut.init = 16'h3aca;
    FD1P3AX block_w2_reg__i1 (.D(n3899[32]), .SP(block_w2_we), .CK(clk_c), 
            .Q(dec_new_block[32])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w2_reg__i1.GSR = "ENABLED";
    LUT4 mux_224_i12_3_lut (.A(dec_new_block[107]), .B(dec_new_block[75]), 
         .C(n6362[1]), .Z(n2752[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam mux_224_i12_3_lut.init = 16'hcaca;
    LUT4 n2763_bdd_4_lut (.A(n2752[21]), .B(n9406), .C(n30146), .D(n25333), 
         .Z(tmp_sboxw[21])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n2763_bdd_4_lut.init = 16'h00ca;
    LUT4 i3_3_lut_4_lut_adj_92 (.A(n33756), .B(n33672), .C(block_new_127__N_1901[105]), 
         .D(block_new_127__N_1901[113]), .Z(n8_adj_7754)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i3_3_lut_4_lut_adj_92.init = 16'h6996;
    LUT4 mux_626_Mux_121_i2_4_lut (.A(new_sboxw[25]), .B(n7_adj_7782), .C(update_type[0]), 
         .D(n8_adj_7687), .Z(n2_adj_7783)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_121_i2_4_lut.init = 16'h3aca;
    LUT4 i27663_3_lut_4_lut (.A(block_new_127__N_1645_c[48]), .B(update_type[0]), 
         .C(n33844), .D(n13076), .Z(n4540[16])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27663_3_lut_4_lut.init = 16'hf808;
    LUT4 i3779_3_lut (.A(dec_new_block[44]), .B(dec_new_block[12]), .C(n6362[3]), 
         .Z(n9388)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam i3779_3_lut.init = 16'hcaca;
    LUT4 mux_626_Mux_0_i2_4_lut (.A(new_sboxw[0]), .B(n29429), .C(update_type[0]), 
         .D(n4_adj_7671), .Z(n2_adj_7784)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_0_i2_4_lut.init = 16'h3aca;
    LUT4 mux_224_i13_3_lut (.A(dec_new_block[108]), .B(dec_new_block[76]), 
         .C(n6362[1]), .Z(n2752[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam mux_224_i13_3_lut.init = 16'hcaca;
    LUT4 mux_626_Mux_2_i2_4_lut (.A(new_sboxw[2]), .B(n5_adj_7785), .C(update_type[0]), 
         .D(n6_adj_7786), .Z(n2_adj_7787)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_2_i2_4_lut.init = 16'h3aca;
    LUT4 i3781_3_lut (.A(dec_new_block[45]), .B(dec_new_block[13]), .C(n6362[3]), 
         .Z(n9390)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam i3781_3_lut.init = 16'hcaca;
    LUT4 mux_626_Mux_6_i2_4_lut (.A(new_sboxw[6]), .B(n7_adj_7788), .C(update_type[0]), 
         .D(n8_adj_7789), .Z(n2_adj_7790)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_6_i2_4_lut.init = 16'h3aca;
    LUT4 mux_224_i14_3_lut (.A(dec_new_block[109]), .B(dec_new_block[77]), 
         .C(n6362[1]), .Z(n2752[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam mux_224_i14_3_lut.init = 16'hcaca;
    LUT4 i3783_3_lut (.A(dec_new_block[46]), .B(dec_new_block[14]), .C(n6362[3]), 
         .Z(n9392)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam i3783_3_lut.init = 16'hcaca;
    LUT4 mux_626_Mux_9_i2_4_lut (.A(new_sboxw[9]), .B(n9_adj_7791), .C(update_type[0]), 
         .D(n10_adj_7792), .Z(n2_adj_7793)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_9_i2_4_lut.init = 16'h3aca;
    FD1P3AY sword_ctr_reg_FSM_i0_i0 (.D(n2689[0]), .SP(sword_ctr_we), .CK(clk_c), 
            .Q(n6362[0]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam sword_ctr_reg_FSM_i0_i0.GSR = "ENABLED";
    LUT4 mux_224_i15_3_lut (.A(dec_new_block[110]), .B(dec_new_block[78]), 
         .C(n6362[1]), .Z(n2752[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam mux_224_i15_3_lut.init = 16'hcaca;
    LUT4 mux_626_Mux_10_i2_4_lut (.A(new_sboxw[10]), .B(n7_adj_7794), .C(update_type[0]), 
         .D(n8_adj_7795), .Z(n2_adj_7796)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_10_i2_4_lut.init = 16'h3aca;
    LUT4 i3785_3_lut (.A(dec_new_block[47]), .B(dec_new_block[15]), .C(n6362[3]), 
         .Z(n9394)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam i3785_3_lut.init = 16'hcaca;
    LUT4 mux_626_Mux_14_i2_4_lut (.A(new_sboxw[14]), .B(n5_adj_7681), .C(update_type[0]), 
         .D(n6_adj_7797), .Z(n2_adj_7798)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_14_i2_4_lut.init = 16'h3aca;
    LUT4 mux_224_i16_3_lut (.A(dec_new_block[111]), .B(dec_new_block[79]), 
         .C(n6362[1]), .Z(n2752[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam mux_224_i16_3_lut.init = 16'hcaca;
    LUT4 i2_2_lut_4_lut_adj_93 (.A(n33583), .B(block_new_127__N_1901[121]), 
         .C(block_new_127__N_1901[114]), .D(n33579), .Z(n6_adj_7786)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i2_2_lut_4_lut_adj_93.init = 16'h6996;
    LUT4 i27511_3_lut_4_lut (.A(block_new_127__N_1645_c[79]), .B(update_type[0]), 
         .C(n33844), .D(n13075), .Z(n4540[15])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27511_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_626_Mux_20_i2_4_lut (.A(new_sboxw[20]), .B(n5_adj_7799), .C(update_type[0]), 
         .D(n6_adj_7800), .Z(n2_adj_7801)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_20_i2_4_lut.init = 16'h3aca;
    LUT4 i3787_3_lut (.A(dec_new_block[48]), .B(dec_new_block[16]), .C(n6362[3]), 
         .Z(n9396)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam i3787_3_lut.init = 16'hcaca;
    LUT4 mux_224_i17_3_lut (.A(dec_new_block[112]), .B(dec_new_block[80]), 
         .C(n6362[1]), .Z(n2752[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam mux_224_i17_3_lut.init = 16'hcaca;
    LUT4 i3789_3_lut (.A(dec_new_block[49]), .B(dec_new_block[17]), .C(n6362[3]), 
         .Z(n9398)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam i3789_3_lut.init = 16'hcaca;
    LUT4 mux_224_i18_3_lut (.A(dec_new_block[113]), .B(dec_new_block[81]), 
         .C(n6362[1]), .Z(n2752[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam mux_224_i18_3_lut.init = 16'hcaca;
    LUT4 i3_3_lut_4_lut_adj_94 (.A(n33697), .B(n33587), .C(n12090), .D(n33779), 
         .Z(n8_adj_7802)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i3_3_lut_4_lut_adj_94.init = 16'h6996;
    LUT4 mux_626_Mux_21_i2_4_lut (.A(new_sboxw[21]), .B(n5_adj_7803), .C(update_type[0]), 
         .D(n6_adj_7804), .Z(n2_adj_7805)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_21_i2_4_lut.init = 16'h3aca;
    LUT4 n2764_bdd_4_lut (.A(n2752[20]), .B(n9404), .C(n30146), .D(n25333), 
         .Z(tmp_sboxw[20])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n2764_bdd_4_lut.init = 16'h00ca;
    LUT4 i3791_3_lut (.A(dec_new_block[50]), .B(dec_new_block[18]), .C(n6362[3]), 
         .Z(n9400)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam i3791_3_lut.init = 16'hcaca;
    LUT4 mux_626_Mux_30_i2_4_lut (.A(new_sboxw[30]), .B(n5_adj_7806), .C(update_type[0]), 
         .D(n6_adj_7807), .Z(n2_adj_7808)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_30_i2_4_lut.init = 16'h3aca;
    LUT4 mux_224_i19_3_lut (.A(dec_new_block[114]), .B(dec_new_block[82]), 
         .C(n6362[1]), .Z(n2752[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam mux_224_i19_3_lut.init = 16'hcaca;
    LUT4 mux_626_Mux_31_i2_4_lut (.A(new_sboxw[31]), .B(n5_adj_7809), .C(update_type[0]), 
         .D(n6_adj_7810), .Z(n2_adj_7811)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_31_i2_4_lut.init = 16'h3aca;
    LUT4 i2_2_lut_4_lut_adj_95 (.A(block_new_127__N_1901[0]), .B(block_new_127__N_1901[14]), 
         .C(n33584), .D(block_new_127__N_1901[23]), .Z(n7_adj_7812)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i2_2_lut_4_lut_adj_95.init = 16'h6996;
    LUT4 i1_2_lut_3_lut_4_lut_adj_96 (.A(block_new_127__N_1901[79]), .B(block_new_127__N_1901[95]), 
         .C(block_new_127__N_1901[71]), .D(n33762), .Z(n4_adj_7813)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_3_lut_4_lut_adj_96.init = 16'h6996;
    LUT4 mux_626_Mux_37_i2_4_lut (.A(new_sboxw[5]), .B(n29273), .C(update_type[0]), 
         .D(n4_adj_7814), .Z(n2_adj_7815)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_37_i2_4_lut.init = 16'h3aca;
    LUT4 i3793_3_lut (.A(dec_new_block[51]), .B(dec_new_block[19]), .C(n6362[3]), 
         .Z(n9402)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam i3793_3_lut.init = 16'hcaca;
    LUT4 i2_2_lut_4_lut_adj_97 (.A(n33524), .B(n648[3]), .C(n873[3]), 
         .D(n29441), .Z(n6_adj_7816)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i2_2_lut_4_lut_adj_97.init = 16'h6996;
    LUT4 mux_626_Mux_38_i2_4_lut (.A(new_sboxw[6]), .B(n9_adj_7817), .C(update_type[0]), 
         .D(n10_adj_7818), .Z(n2_adj_7819)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_38_i2_4_lut.init = 16'h3aca;
    LUT4 mux_224_i20_3_lut (.A(dec_new_block[115]), .B(dec_new_block[83]), 
         .C(n6362[1]), .Z(n2752[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam mux_224_i20_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut_adj_98 (.A(block_new_127__N_1901[0]), .B(block_new_127__N_1901[14]), 
         .C(n33584), .D(n33828), .Z(n4_adj_7820)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_4_lut_adj_98.init = 16'h6996;
    LUT4 i2_2_lut_4_lut_adj_99 (.A(n33698), .B(block_new_127__N_1901[45]), 
         .C(n4770[4]), .D(n33671), .Z(n6_adj_7775)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i2_2_lut_4_lut_adj_99.init = 16'h6996;
    LUT4 mux_626_Mux_41_i2_4_lut (.A(new_sboxw[9]), .B(n5_adj_7821), .C(update_type[0]), 
         .D(n6_adj_7822), .Z(n2_adj_7823)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_41_i2_4_lut.init = 16'h3aca;
    LUT4 i3795_3_lut (.A(dec_new_block[52]), .B(dec_new_block[20]), .C(n6362[3]), 
         .Z(n9404)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam i3795_3_lut.init = 16'hcaca;
    LUT4 mux_224_i21_3_lut (.A(dec_new_block[116]), .B(dec_new_block[84]), 
         .C(n6362[1]), .Z(n2752[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam mux_224_i21_3_lut.init = 16'hcaca;
    LUT4 mux_626_Mux_42_i2_4_lut (.A(new_sboxw[10]), .B(n7_adj_7677), .C(update_type[0]), 
         .D(n8_adj_7824), .Z(n2_adj_7825)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_42_i2_4_lut.init = 16'h3aca;
    LUT4 i3797_3_lut (.A(dec_new_block[53]), .B(dec_new_block[21]), .C(n6362[3]), 
         .Z(n9406)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam i3797_3_lut.init = 16'hcaca;
    LUT4 mux_224_i22_3_lut (.A(dec_new_block[117]), .B(dec_new_block[85]), 
         .C(n6362[1]), .Z(n2752[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam mux_224_i22_3_lut.init = 16'hcaca;
    LUT4 mux_626_Mux_47_i2_4_lut (.A(new_sboxw[15]), .B(n33769), .C(update_type[0]), 
         .D(n4_adj_7826), .Z(n2_adj_7827)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_47_i2_4_lut.init = 16'h3aca;
    LUT4 i3799_3_lut (.A(dec_new_block[54]), .B(dec_new_block[22]), .C(n6362[3]), 
         .Z(n9408)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam i3799_3_lut.init = 16'hcaca;
    LUT4 mux_626_Mux_60_i2_4_lut (.A(new_sboxw[28]), .B(n33520), .C(update_type[0]), 
         .D(n4_adj_7672), .Z(n2_adj_7828)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_60_i2_4_lut.init = 16'h3aca;
    LUT4 mux_224_i23_3_lut (.A(dec_new_block[118]), .B(dec_new_block[86]), 
         .C(n6362[1]), .Z(n2752[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam mux_224_i23_3_lut.init = 16'hcaca;
    LUT4 i3_3_lut_4_lut_adj_100 (.A(block_new_127__N_1901[53]), .B(n33586), 
         .C(n33812), .D(n33799), .Z(n8_adj_7829)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i3_3_lut_4_lut_adj_100.init = 16'h6996;
    LUT4 mux_626_Mux_66_i2_4_lut (.A(new_sboxw[2]), .B(n9_adj_7830), .C(update_type[0]), 
         .D(n10_adj_7831), .Z(n2_adj_7832)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_66_i2_4_lut.init = 16'h3aca;
    FD1S3AY ready_reg_830 (.D(n6431), .CK(clk_c), .Q(dec_ready));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam ready_reg_830.GSR = "ENABLED";
    LUT4 i3801_3_lut (.A(dec_new_block[55]), .B(dec_new_block[23]), .C(n6362[3]), 
         .Z(n9410)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam i3801_3_lut.init = 16'hcaca;
    LUT4 mux_224_i24_3_lut (.A(dec_new_block[119]), .B(dec_new_block[87]), 
         .C(n6362[1]), .Z(n2752[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam mux_224_i24_3_lut.init = 16'hcaca;
    LUT4 n2765_bdd_4_lut (.A(n2752[19]), .B(n9402), .C(n30146), .D(n25333), 
         .Z(tmp_sboxw[19])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n2765_bdd_4_lut.init = 16'h00ca;
    LUT4 mux_626_Mux_67_i2_4_lut (.A(new_sboxw[3]), .B(n9_adj_7833), .C(update_type[0]), 
         .D(n10_adj_7834), .Z(n2_adj_7835)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_67_i2_4_lut.init = 16'h3aca;
    LUT4 i3803_3_lut (.A(dec_new_block[56]), .B(dec_new_block[24]), .C(n6362[3]), 
         .Z(n9412)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam i3803_3_lut.init = 16'hcaca;
    LUT4 mux_224_i25_3_lut (.A(dec_new_block[120]), .B(dec_new_block[88]), 
         .C(n6362[1]), .Z(n2752[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam mux_224_i25_3_lut.init = 16'hcaca;
    LUT4 mux_626_Mux_68_i2_4_lut (.A(new_sboxw[4]), .B(n5_adj_7836), .C(update_type[0]), 
         .D(n6_adj_7837), .Z(n2_adj_7838)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_68_i2_4_lut.init = 16'h3aca;
    LUT4 i3805_3_lut (.A(dec_new_block[57]), .B(dec_new_block[25]), .C(n6362[3]), 
         .Z(n9414)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam i3805_3_lut.init = 16'hcaca;
    LUT4 mux_224_i26_3_lut (.A(dec_new_block[121]), .B(dec_new_block[89]), 
         .C(n6362[1]), .Z(n2752[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam mux_224_i26_3_lut.init = 16'hcaca;
    LUT4 mux_626_Mux_74_i2_4_lut (.A(new_sboxw[10]), .B(n28882), .C(update_type[0]), 
         .D(n4_adj_7839), .Z(n2_adj_7840)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_74_i2_4_lut.init = 16'h3aca;
    LUT4 mux_626_Mux_77_i2_4_lut (.A(new_sboxw[13]), .B(n33519), .C(update_type[0]), 
         .D(n4_adj_7841), .Z(n2_adj_7842)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_77_i2_4_lut.init = 16'h3aca;
    LUT4 i3807_3_lut (.A(dec_new_block[58]), .B(dec_new_block[26]), .C(n6362[3]), 
         .Z(n9416)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam i3807_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_101 (.A(n33699), .B(n33706), .C(n33800), 
         .D(block_new_127__N_1901[53]), .Z(n4_adj_7843)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_3_lut_4_lut_adj_101.init = 16'h6996;
    FD1P3AX dec_ctrl_reg_FSM_i0_i0 (.D(n149), .SP(dec_ctrl_we), .CK(clk_c), 
            .Q(n6363[0]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(462[7] 518[14])
    defparam dec_ctrl_reg_FSM_i0_i0.GSR = "ENABLED";
    LUT4 mux_626_Mux_78_i2_4_lut (.A(new_sboxw[14]), .B(n5_adj_7844), .C(update_type[0]), 
         .D(n6_adj_7845), .Z(n2_adj_7846)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_78_i2_4_lut.init = 16'h3aca;
    LUT4 mux_224_i27_3_lut (.A(dec_new_block[122]), .B(dec_new_block[90]), 
         .C(n6362[1]), .Z(n2752[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam mux_224_i27_3_lut.init = 16'hcaca;
    LUT4 mux_626_Mux_81_i2_4_lut (.A(new_sboxw[17]), .B(n7_adj_7847), .C(update_type[0]), 
         .D(n8_adj_7848), .Z(n2_adj_7849)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_81_i2_4_lut.init = 16'h3aca;
    LUT4 mux_626_Mux_88_i2_4_lut (.A(new_sboxw[24]), .B(n7_adj_7850), .C(update_type[0]), 
         .D(n8_adj_7851), .Z(n2_adj_7852)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_88_i2_4_lut.init = 16'h3aca;
    LUT4 i3809_3_lut (.A(dec_new_block[59]), .B(dec_new_block[27]), .C(n6362[3]), 
         .Z(n9418)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam i3809_3_lut.init = 16'hcaca;
    LUT4 mux_224_i28_3_lut (.A(dec_new_block[123]), .B(dec_new_block[91]), 
         .C(n6362[1]), .Z(n2752[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam mux_224_i28_3_lut.init = 16'hcaca;
    LUT4 mux_626_Mux_90_i2_4_lut (.A(new_sboxw[26]), .B(n5_adj_7853), .C(update_type[0]), 
         .D(n6_adj_7854), .Z(n2_adj_7855)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_90_i2_4_lut.init = 16'h3aca;
    LUT4 new_block_127__I_0_i123_2_lut (.A(dec_new_block[122]), .B(round_key[122]), 
         .Z(block_new_127__N_1901[122])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i123_2_lut.init = 16'h6666;
    LUT4 i3811_3_lut (.A(dec_new_block[60]), .B(dec_new_block[28]), .C(n6362[3]), 
         .Z(n9420)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam i3811_3_lut.init = 16'hcaca;
    LUT4 mux_626_Mux_94_i2_4_lut (.A(new_sboxw[30]), .B(n5_adj_7856), .C(update_type[0]), 
         .D(n6_adj_7679), .Z(n2_adj_7857)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_94_i2_4_lut.init = 16'h3aca;
    LUT4 mux_224_i29_3_lut (.A(dec_new_block[124]), .B(dec_new_block[92]), 
         .C(n6362[1]), .Z(n2752[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam mux_224_i29_3_lut.init = 16'hcaca;
    LUT4 i27589_3_lut_4_lut (.A(block_new_127__N_1645_c[78]), .B(update_type[0]), 
         .C(n33844), .D(n13074), .Z(n4540[14])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27589_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_626_Mux_95_i2_4_lut (.A(new_sboxw[31]), .B(n29244), .C(update_type[0]), 
         .D(n4_adj_7858), .Z(n2_adj_7859)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_95_i2_4_lut.init = 16'h3aca;
    LUT4 i3813_3_lut (.A(dec_new_block[61]), .B(dec_new_block[29]), .C(n6362[3]), 
         .Z(n9422)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam i3813_3_lut.init = 16'hcaca;
    LUT4 mux_224_i30_3_lut (.A(dec_new_block[125]), .B(dec_new_block[93]), 
         .C(n6362[1]), .Z(n2752[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam mux_224_i30_3_lut.init = 16'hcaca;
    LUT4 mux_626_Mux_102_i2_4_lut (.A(new_sboxw[6]), .B(n7_adj_7860), .C(update_type[0]), 
         .D(n8_adj_7682), .Z(n2_adj_7861)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_102_i2_4_lut.init = 16'h3aca;
    LUT4 i27653_3_lut_4_lut (.A(block_new_127__N_1645_c[127]), .B(update_type[0]), 
         .C(n33844), .D(n13187), .Z(n4540[127])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27653_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_626_Mux_109_i2_4_lut (.A(new_sboxw[13]), .B(n7_adj_7862), .C(update_type[0]), 
         .D(n8_adj_7684), .Z(n2_adj_7863)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_109_i2_4_lut.init = 16'h3aca;
    LUT4 i27651_3_lut_4_lut (.A(block_new_127__N_1645_c[126]), .B(update_type[0]), 
         .C(n33844), .D(n13186), .Z(n4540[126])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27651_3_lut_4_lut.init = 16'hf808;
    LUT4 i3815_3_lut (.A(dec_new_block[62]), .B(dec_new_block[30]), .C(n6362[3]), 
         .Z(n9424)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam i3815_3_lut.init = 16'hcaca;
    LUT4 mux_626_Mux_111_i2_4_lut (.A(new_sboxw[15]), .B(n5_adj_7864), .C(update_type[0]), 
         .D(n6_adj_7689), .Z(n2_adj_7865)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_111_i2_4_lut.init = 16'h3aca;
    LUT4 mux_224_i31_3_lut (.A(dec_new_block[126]), .B(dec_new_block[94]), 
         .C(n6362[1]), .Z(n2752[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam mux_224_i31_3_lut.init = 16'hcaca;
    LUT4 mux_626_Mux_113_i2_4_lut (.A(new_sboxw[17]), .B(n9_adj_7866), .C(update_type[0]), 
         .D(n10_adj_7867), .Z(n2_adj_7868)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_113_i2_4_lut.init = 16'h3aca;
    LUT4 i3817_3_lut (.A(dec_new_block[63]), .B(dec_new_block[31]), .C(n6362[3]), 
         .Z(n9426)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam i3817_3_lut.init = 16'hcaca;
    LUT4 i27509_3_lut_4_lut (.A(block_new_127__N_1645_c[77]), .B(update_type[0]), 
         .C(n33844), .D(n13073), .Z(n4540[13])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27509_3_lut_4_lut.init = 16'hf808;
    LUT4 i27661_3_lut_4_lut (.A(\block_new_127__N_1645[76] ), .B(update_type[0]), 
         .C(n33844), .D(n13072), .Z(n4540[12])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27661_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_224_i32_3_lut (.A(dec_new_block[127]), .B(dec_new_block[95]), 
         .C(n6362[1]), .Z(n2752[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam mux_224_i32_3_lut.init = 16'hcaca;
    LUT4 mux_626_Mux_116_i2_4_lut (.A(new_sboxw[20]), .B(n29291), .C(update_type[0]), 
         .D(n4_adj_7869), .Z(n2_adj_7870)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_116_i2_4_lut.init = 16'h3aca;
    LUT4 i2_2_lut_4_lut_adj_102 (.A(n33804), .B(block_new_127__N_1901[78]), 
         .C(n33590), .D(block_new_127__N_1901[72]), .Z(n7_adj_7871)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i2_2_lut_4_lut_adj_102.init = 16'h6996;
    LUT4 mux_626_Mux_117_i2_4_lut (.A(new_sboxw[21]), .B(n29273), .C(update_type[0]), 
         .D(n4_adj_7872), .Z(n2_adj_7873)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_117_i2_4_lut.init = 16'h3aca;
    LUT4 i27797_3_lut_4_lut (.A(\block_new_127__N_1645[125] ), .B(update_type[0]), 
         .C(n33844), .D(n13185), .Z(n4540[125])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27797_3_lut_4_lut.init = 16'hf808;
    LUT4 i27649_3_lut_4_lut (.A(block_new_127__N_1645_c[124]), .B(update_type[0]), 
         .C(n33844), .D(n13184), .Z(n4540[124])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27649_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_626_Mux_118_i2_4_lut (.A(new_sboxw[22]), .B(n7_adj_7874), .C(update_type[0]), 
         .D(n8_adj_7875), .Z(n2_adj_7876)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_118_i2_4_lut.init = 16'h3aca;
    LUT4 new_block_127__I_0_i1_2_lut (.A(dec_new_block[0]), .B(round_key[0]), 
         .Z(block_new_127__N_1901[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i1_2_lut.init = 16'h6666;
    LUT4 i9301_3_lut (.A(dec_round_nr_c[1]), .B(dec_round_nr_c[2]), .C(dec_round_nr[0]), 
         .Z(n14912)) /* synthesis lut_function=(A (B)+!A (B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(99[18:30])
    defparam i9301_3_lut.init = 16'hc9c9;
    LUT4 i27795_3_lut_4_lut (.A(\block_new_127__N_1645[123] ), .B(update_type[0]), 
         .C(n33844), .D(n13183), .Z(n4540[123])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27795_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_626_Mux_122_i2_4_lut (.A(new_sboxw[26]), .B(n7_adj_7877), .C(update_type[0]), 
         .D(n8_adj_7878), .Z(n2_adj_7879)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_122_i2_4_lut.init = 16'h3aca;
    LUT4 i27853_4_lut (.A(\key_mem_ctrl.num_rounds[2] ), .B(encdec_reg), 
         .C(n149), .D(\aes_core_ctrl_new_1__N_858[1] ), .Z(n30080)) /* synthesis lut_function=(!(A (B+!(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_key_mem.v(366[19:29])
    defparam i27853_4_lut.init = 16'h7555;
    LUT4 i1_2_lut (.A(\aes_core_ctrl_new_1__N_858[1] ), .B(encdec_reg), 
         .Z(n110)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(96[7:17])
    defparam i1_2_lut.init = 16'h2222;
    LUT4 i9631_3_lut (.A(dec_round_nr_c[3]), .B(\enc_round_nr[3] ), .C(encdec_reg), 
         .Z(\muxed_round_nr[3] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(96[7:17])
    defparam i9631_3_lut.init = 16'hcaca;
    LUT4 i9397_3_lut (.A(dec_round_nr_c[2]), .B(\enc_round_nr[2] ), .C(encdec_reg), 
         .Z(\muxed_round_nr[2] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(96[7:17])
    defparam i9397_3_lut.init = 16'hcaca;
    LUT4 i27647_3_lut_4_lut (.A(block_new_127__N_1645_c[122]), .B(update_type[0]), 
         .C(n33844), .D(n13182), .Z(n4540[122])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27647_3_lut_4_lut.init = 16'hf808;
    LUT4 i27577_3_lut_4_lut (.A(\block_new_127__N_1645[121] ), .B(update_type[0]), 
         .C(n33844), .D(n13181), .Z(n4540[121])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27577_3_lut_4_lut.init = 16'hf808;
    LUT4 i27575_3_lut_4_lut (.A(block_new_127__N_1645_c[120]), .B(update_type[0]), 
         .C(n33844), .D(n13180), .Z(n4540[120])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27575_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_626_Mux_124_i2_4_lut (.A(new_sboxw[28]), .B(n7_adj_7880), .C(update_type[0]), 
         .D(n8_adj_7881), .Z(n2_adj_7882)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_124_i2_4_lut.init = 16'h3aca;
    LUT4 mux_626_Mux_126_i2_4_lut (.A(new_sboxw[30]), .B(n7_adj_7883), .C(update_type[0]), 
         .D(n8_adj_7718), .Z(n2_adj_7884)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_126_i2_4_lut.init = 16'h3aca;
    LUT4 mux_626_Mux_127_i2_4_lut (.A(new_sboxw[31]), .B(n5_adj_7885), .C(update_type[0]), 
         .D(n6_adj_7886), .Z(n2_adj_7887)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_127_i2_4_lut.init = 16'h3aca;
    LUT4 i27249_3_lut_4_lut (.A(block_new_127__N_1645_c[23]), .B(update_type[0]), 
         .C(n33844), .D(n13179), .Z(n4540[119])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27249_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_626_Mux_3_i2_4_lut (.A(new_sboxw[3]), .B(n7_adj_7888), .C(update_type[0]), 
         .D(n8_adj_7889), .Z(n2_adj_7890)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_3_i2_4_lut.init = 16'h3aca;
    LUT4 i27645_3_lut_4_lut (.A(block_new_127__N_1645_c[22]), .B(update_type[0]), 
         .C(n33844), .D(n13178), .Z(n4540[118])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27645_3_lut_4_lut.init = 16'hf808;
    LUT4 i27643_3_lut_4_lut (.A(\block_new_127__N_1645[21] ), .B(update_type[0]), 
         .C(n33844), .D(n13177), .Z(n4540[117])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27643_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_626_Mux_4_i2_4_lut (.A(new_sboxw[4]), .B(n29462), .C(update_type[0]), 
         .D(n4_adj_7891), .Z(n2_adj_7892)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_4_i2_4_lut.init = 16'h3aca;
    LUT4 mux_626_Mux_8_i2_4_lut (.A(new_sboxw[8]), .B(n33521), .C(update_type[0]), 
         .D(n4_adj_7893), .Z(n2_adj_7894)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_8_i2_4_lut.init = 16'h3aca;
    LUT4 i27641_3_lut_4_lut (.A(\block_new_127__N_1645[20] ), .B(update_type[0]), 
         .C(n33844), .D(n13176), .Z(n4540[116])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27641_3_lut_4_lut.init = 16'hf808;
    LUT4 i27751_3_lut_4_lut (.A(\block_new_127__N_1645[19] ), .B(update_type[0]), 
         .C(n33844), .D(n13175), .Z(n4540[115])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27751_3_lut_4_lut.init = 16'hf808;
    LUT4 i27247_3_lut_4_lut (.A(block_new_127__N_1645_c[18]), .B(update_type[0]), 
         .C(n33844), .D(n13174), .Z(n4540[114])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27247_3_lut_4_lut.init = 16'hf808;
    LUT4 n2766_bdd_4_lut (.A(n2752[18]), .B(n9400), .C(n30146), .D(n25333), 
         .Z(tmp_sboxw[18])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n2766_bdd_4_lut.init = 16'h00ca;
    LUT4 block_127__I_0_i125_2_lut (.A(\block_reg[0] [28]), .B(round_key[124]), 
         .Z(block_new_127__N_1645_c[124])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i125_2_lut.init = 16'h6666;
    LUT4 i27639_3_lut_4_lut (.A(\block_new_127__N_1645[17] ), .B(update_type[0]), 
         .C(n33844), .D(n13173), .Z(n4540[113])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27639_3_lut_4_lut.init = 16'hf808;
    LUT4 i27573_3_lut_4_lut (.A(block_new_127__N_1645_c[16]), .B(update_type[0]), 
         .C(n33844), .D(n13172), .Z(n4540[112])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27573_3_lut_4_lut.init = 16'hf808;
    LUT4 i27637_3_lut_4_lut (.A(block_new_127__N_1645_c[47]), .B(update_type[0]), 
         .C(n33844), .D(n13171), .Z(n4540[111])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27637_3_lut_4_lut.init = 16'hf808;
    LUT4 i27571_3_lut_4_lut (.A(block_new_127__N_1645_c[46]), .B(update_type[0]), 
         .C(n33844), .D(n13170), .Z(n4540[110])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27571_3_lut_4_lut.init = 16'hf808;
    LUT4 i27635_3_lut_4_lut (.A(block_new_127__N_1645_c[45]), .B(update_type[0]), 
         .C(n33844), .D(n13169), .Z(n4540[109])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27635_3_lut_4_lut.init = 16'hf808;
    LUT4 i27709_3_lut_4_lut (.A(\block_new_127__N_1645[44] ), .B(update_type[0]), 
         .C(n33844), .D(n13168), .Z(n4540[108])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27709_3_lut_4_lut.init = 16'hf808;
    LUT4 i27749_3_lut_4_lut (.A(\block_new_127__N_1645[43] ), .B(update_type[0]), 
         .C(n33844), .D(n13167), .Z(n4540[107])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27749_3_lut_4_lut.init = 16'hf808;
    LUT4 i27569_3_lut_4_lut (.A(block_new_127__N_1645_c[42]), .B(update_type[0]), 
         .C(n33844), .D(n13166), .Z(n4540[106])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27569_3_lut_4_lut.init = 16'hf808;
    LUT4 i27747_3_lut_4_lut (.A(\block_new_127__N_1645[41] ), .B(update_type[0]), 
         .C(n33844), .D(n13165), .Z(n4540[105])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27747_3_lut_4_lut.init = 16'hf808;
    LUT4 i27567_3_lut_4_lut (.A(block_new_127__N_1645_c[40]), .B(update_type[0]), 
         .C(n33844), .D(n13164), .Z(n4540[104])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27567_3_lut_4_lut.init = 16'hf808;
    LUT4 i27565_3_lut_4_lut (.A(\block_new_127__N_1645[71] ), .B(update_type[0]), 
         .C(n33844), .D(n13163), .Z(n4540[103])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27565_3_lut_4_lut.init = 16'hf808;
    LUT4 i27633_3_lut_4_lut (.A(\block_new_127__N_1645[70] ), .B(update_type[0]), 
         .C(n33844), .D(n13162), .Z(n4540[102])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27633_3_lut_4_lut.init = 16'hf808;
    LUT4 i27707_3_lut_4_lut (.A(\block_new_127__N_1645[69] ), .B(update_type[0]), 
         .C(n33844), .D(n13161), .Z(n4540[101])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27707_3_lut_4_lut.init = 16'hf808;
    LUT4 i27705_3_lut_4_lut (.A(\block_new_127__N_1645[68] ), .B(update_type[0]), 
         .C(n33844), .D(n13160), .Z(n4540[100])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27705_3_lut_4_lut.init = 16'hf808;
    LUT4 i27703_3_lut_4_lut (.A(\block_new_127__N_1645[67] ), .B(update_type[0]), 
         .C(n33844), .D(n13159), .Z(n4540[99])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27703_3_lut_4_lut.init = 16'hf808;
    LUT4 i1_2_lut_adj_103 (.A(n6363[1]), .B(n6362[3]), .Z(n149)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam i1_2_lut_adj_103.init = 16'h8888;
    LUT4 i27563_3_lut_4_lut (.A(block_new_127__N_1645_c[66]), .B(update_type[0]), 
         .C(n33844), .D(n13158), .Z(n4540[98])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27563_3_lut_4_lut.init = 16'hf808;
    LUT4 i27561_3_lut_4_lut (.A(\block_new_127__N_1645[65] ), .B(update_type[0]), 
         .C(n33844), .D(n13157), .Z(n4540[97])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27561_3_lut_4_lut.init = 16'hf808;
    LUT4 i27559_3_lut_4_lut (.A(\block_new_127__N_1645[64] ), .B(update_type[0]), 
         .C(n33844), .D(n13156), .Z(n4540[96])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27559_3_lut_4_lut.init = 16'hf808;
    LUT4 i27631_3_lut_4_lut (.A(block_new_127__N_1645_c[95]), .B(update_type[0]), 
         .C(n33844), .D(n13155), .Z(n4540[95])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27631_3_lut_4_lut.init = 16'hf808;
    LUT4 i27629_3_lut_4_lut (.A(block_new_127__N_1645_c[94]), .B(update_type[0]), 
         .C(n33844), .D(n13154), .Z(n4540[94])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27629_3_lut_4_lut.init = 16'hf808;
    LUT4 i27701_3_lut_4_lut (.A(block_new_127__N_1645_c[93]), .B(update_type[0]), 
         .C(n33844), .D(n13153), .Z(n4540[93])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27701_3_lut_4_lut.init = 16'hf808;
    LUT4 i27699_3_lut_4_lut (.A(\block_new_127__N_1645[92] ), .B(update_type[0]), 
         .C(n33844), .D(n13152), .Z(n4540[92])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27699_3_lut_4_lut.init = 16'hf808;
    LUT4 i27745_3_lut_4_lut (.A(\block_new_127__N_1645[91] ), .B(update_type[0]), 
         .C(n33844), .D(n13151), .Z(n4540[91])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27745_3_lut_4_lut.init = 16'hf808;
    LUT4 i27627_3_lut_4_lut (.A(block_new_127__N_1645_c[90]), .B(update_type[0]), 
         .C(n33844), .D(n13150), .Z(n4540[90])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27627_3_lut_4_lut.init = 16'hf808;
    LUT4 i27557_3_lut_4_lut (.A(\block_new_127__N_1645[89] ), .B(update_type[0]), 
         .C(n33844), .D(n13149), .Z(n4540[89])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27557_3_lut_4_lut.init = 16'hf808;
    LUT4 i27625_3_lut_4_lut (.A(block_new_127__N_1645_c[88]), .B(update_type[0]), 
         .C(n33844), .D(n13148), .Z(n4540[88])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27625_3_lut_4_lut.init = 16'hf808;
    LUT4 i27245_3_lut_4_lut (.A(\block_new_127__N_1645[119] ), .B(update_type[0]), 
         .C(n33844), .D(n13147), .Z(n4540[87])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27245_3_lut_4_lut.init = 16'hf808;
    LUT4 i27555_3_lut_4_lut (.A(\block_new_127__N_1645[118] ), .B(update_type[0]), 
         .C(n33844), .D(n13146), .Z(n4540[86])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27555_3_lut_4_lut.init = 16'hf808;
    LUT4 i27743_3_lut_4_lut (.A(block_new_127__N_1645_c[117]), .B(update_type[0]), 
         .C(n33844), .D(n13145), .Z(n4540[85])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27743_3_lut_4_lut.init = 16'hf808;
    LUT4 i27697_3_lut_4_lut (.A(\block_new_127__N_1645[116] ), .B(update_type[0]), 
         .C(n33844), .D(n13144), .Z(n4540[84])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27697_3_lut_4_lut.init = 16'hf808;
    LUT4 i27793_3_lut_4_lut (.A(\block_new_127__N_1645[115] ), .B(update_type[0]), 
         .C(n33844), .D(n13143), .Z(n4540[83])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27793_3_lut_4_lut.init = 16'hf808;
    LUT4 i27553_3_lut_4_lut (.A(\block_new_127__N_1645[114] ), .B(update_type[0]), 
         .C(n33844), .D(n13142), .Z(n4540[82])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27553_3_lut_4_lut.init = 16'hf808;
    LUT4 i27623_3_lut_4_lut (.A(\block_new_127__N_1645[113] ), .B(update_type[0]), 
         .C(n33844), .D(n13141), .Z(n4540[81])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27623_3_lut_4_lut.init = 16'hf808;
    LUT4 i27551_3_lut_4_lut (.A(block_new_127__N_1645_c[112]), .B(update_type[0]), 
         .C(n33844), .D(n13140), .Z(n4540[80])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27551_3_lut_4_lut.init = 16'hf808;
    LUT4 i27549_3_lut_4_lut (.A(block_new_127__N_1645_c[15]), .B(update_type[0]), 
         .C(n33844), .D(n13139), .Z(n4540[79])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27549_3_lut_4_lut.init = 16'hf808;
    LUT4 i27621_3_lut_4_lut (.A(\block_new_127__N_1645[14] ), .B(update_type[0]), 
         .C(n33844), .D(n13138), .Z(n4540[78])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27621_3_lut_4_lut.init = 16'hf808;
    LUT4 n2767_bdd_4_lut (.A(n2752[17]), .B(n9398), .C(n30146), .D(n25333), 
         .Z(tmp_sboxw[17])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n2767_bdd_4_lut.init = 16'h00ca;
    LUT4 i27619_3_lut_4_lut (.A(block_new_127__N_1645_c[13]), .B(update_type[0]), 
         .C(n33844), .D(n13137), .Z(n4540[77])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27619_3_lut_4_lut.init = 16'hf808;
    LUT4 block_127__I_0_i124_2_lut (.A(\block_reg[0] [27]), .B(round_key[123]), 
         .Z(\block_new_127__N_1645[123] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i124_2_lut.init = 16'h6666;
    LUT4 i27695_3_lut_4_lut (.A(\block_new_127__N_1645[12] ), .B(update_type[0]), 
         .C(n33844), .D(n13136), .Z(n4540[76])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27695_3_lut_4_lut.init = 16'hf808;
    LUT4 i2_2_lut_4_lut_adj_104 (.A(n33674), .B(block_new_127__N_1901[23]), 
         .C(n33782), .D(block_new_127__N_1901[22]), .Z(n6_adj_7810)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i2_2_lut_4_lut_adj_104.init = 16'h6996;
    LUT4 i27791_3_lut_4_lut (.A(block_new_127__N_1645_c[11]), .B(update_type[0]), 
         .C(n33844), .D(n13135), .Z(n4540[75])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27791_3_lut_4_lut.init = 16'hf808;
    LUT4 i27617_3_lut_4_lut (.A(\block_new_127__N_1645[10] ), .B(update_type[0]), 
         .C(n33844), .D(n13134), .Z(n4540[74])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27617_3_lut_4_lut.init = 16'hf808;
    LUT4 n2768_bdd_4_lut (.A(n2752[16]), .B(n9396), .C(n30146), .D(n25333), 
         .Z(tmp_sboxw[16])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n2768_bdd_4_lut.init = 16'h00ca;
    LUT4 i27547_3_lut_4_lut (.A(block_new_127__N_1645_c[9]), .B(update_type[0]), 
         .C(n33844), .D(n13133), .Z(n4540[73])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27547_3_lut_4_lut.init = 16'hf808;
    LUT4 i2_2_lut_4_lut_adj_105 (.A(n33679), .B(block_new_127__N_1901[127]), 
         .C(n33766), .D(n33758), .Z(n6_adj_7822)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i2_2_lut_4_lut_adj_105.init = 16'h6996;
    LUT4 i27243_3_lut_4_lut (.A(block_new_127__N_1645_c[8]), .B(update_type[0]), 
         .C(n33844), .D(n13132), .Z(n4540[72])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27243_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_626_Mux_12_i2_4_lut (.A(new_sboxw[12]), .B(n5_adj_7896), .C(update_type[0]), 
         .D(n6_adj_7897), .Z(n2_adj_7898)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_12_i2_4_lut.init = 16'h3aca;
    LUT4 mux_626_Mux_16_i2_4_lut (.A(new_sboxw[16]), .B(n33693), .C(update_type[0]), 
         .D(n4_adj_7899), .Z(n2_adj_7900)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_16_i2_4_lut.init = 16'h3aca;
    LUT4 mux_626_Mux_19_i2_4_lut (.A(new_sboxw[19]), .B(n5_adj_7901), .C(update_type[0]), 
         .D(n6_adj_7902), .Z(n2_adj_7903)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_19_i2_4_lut.init = 16'h3aca;
    LUT4 mux_626_Mux_24_i2_4_lut (.A(new_sboxw[24]), .B(n33773), .C(update_type[0]), 
         .D(n4_adj_7820), .Z(n2_adj_7904)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_24_i2_4_lut.init = 16'h3aca;
    LUT4 mux_626_Mux_26_i2_4_lut (.A(new_sboxw[26]), .B(n33777), .C(update_type[0]), 
         .D(n4_adj_7905), .Z(n2_adj_7906)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_26_i2_4_lut.init = 16'h3aca;
    LUT4 i1_2_lut_4_lut_adj_106 (.A(n29444), .B(block_new_127__N_1901[124]), 
         .C(block_new_127__N_1901[109]), .D(n33808), .Z(n5_adj_7907)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_4_lut_adj_106.init = 16'h6996;
    LUT4 i2_2_lut_3_lut_4_lut_adj_107 (.A(block_new_127__N_1901[109]), .B(block_new_127__N_1901[126]), 
         .C(block_new_127__N_1901[102]), .D(block_new_127__N_1901[110]), 
         .Z(n7_adj_7756)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i2_2_lut_3_lut_4_lut_adj_107.init = 16'h6996;
    LUT4 mux_626_Mux_28_i2_4_lut (.A(new_sboxw[28]), .B(n5_adj_7908), .C(update_type[0]), 
         .D(n6_adj_7909), .Z(n2_adj_7910)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_28_i2_4_lut.init = 16'h3aca;
    LUT4 i1_2_lut_4_lut_adj_108 (.A(n29444), .B(block_new_127__N_1901[124]), 
         .C(block_new_127__N_1901[109]), .D(n33807), .Z(n29462)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_4_lut_adj_108.init = 16'h6996;
    LUT4 mux_626_Mux_29_i2_4_lut (.A(new_sboxw[29]), .B(n7_adj_7911), .C(update_type[0]), 
         .D(n8_adj_7802), .Z(n2_adj_7912)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_29_i2_4_lut.init = 16'h3aca;
    LUT4 mux_626_Mux_33_i2_4_lut (.A(new_sboxw[1]), .B(n7_adj_7812), .C(update_type[0]), 
         .D(n8_adj_7913), .Z(n2_adj_7914)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_33_i2_4_lut.init = 16'h3aca;
    LUT4 mux_626_Mux_35_i2_4_lut (.A(new_sboxw[3]), .B(n5_adj_7915), .C(update_type[0]), 
         .D(n6_adj_7916), .Z(n2_adj_7917)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_35_i2_4_lut.init = 16'h3aca;
    LUT4 mux_626_Mux_36_i2_4_lut (.A(new_sboxw[4]), .B(n5_adj_7918), .C(update_type[0]), 
         .D(n6_adj_7919), .Z(n2_adj_7920)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_36_i2_4_lut.init = 16'h3aca;
    LUT4 mux_626_Mux_44_i2_4_lut (.A(new_sboxw[12]), .B(n29462), .C(update_type[0]), 
         .D(n4_adj_7921), .Z(n2_adj_7922)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_44_i2_4_lut.init = 16'h3aca;
    LUT4 i2_2_lut_3_lut_4_lut_adj_109 (.A(n33790), .B(n33715), .C(n33701), 
         .D(n33837), .Z(n6_adj_7923)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i2_2_lut_3_lut_4_lut_adj_109.init = 16'h6996;
    LUT4 i2_2_lut_3_lut_4_lut_adj_110 (.A(block_new_127__N_1901[109]), .B(block_new_127__N_1901[126]), 
         .C(block_new_127__N_1901[103]), .D(block_new_127__N_1901[110]), 
         .Z(n7_adj_7716)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i2_2_lut_3_lut_4_lut_adj_110.init = 16'h6996;
    LUT4 mux_626_Mux_45_i2_4_lut (.A(new_sboxw[13]), .B(n5_adj_7924), .C(update_type[0]), 
         .D(n6_adj_7923), .Z(n2_adj_7925)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_45_i2_4_lut.init = 16'h3aca;
    LUT4 mux_626_Mux_52_i2_4_lut (.A(new_sboxw[20]), .B(n5_adj_7926), .C(update_type[0]), 
         .D(n6_adj_7927), .Z(n2_adj_7928)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_52_i2_4_lut.init = 16'h3aca;
    LUT4 mux_626_Mux_53_i2_4_lut (.A(new_sboxw[21]), .B(n5), .C(update_type[0]), 
         .D(n6_adj_7929), .Z(n2_adj_7930)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_53_i2_4_lut.init = 16'h3aca;
    LUT4 mux_626_Mux_61_i2_4_lut (.A(new_sboxw[29]), .B(n33585), .C(update_type[0]), 
         .D(n4_adj_7843), .Z(n2_adj_7931)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_61_i2_4_lut.init = 16'h3aca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_111 (.A(n33790), .B(n33715), .C(block_new_127__N_1901[116]), 
         .D(n33837), .Z(n4_adj_7891)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_3_lut_4_lut_adj_111.init = 16'h6996;
    LUT4 mux_626_Mux_64_i2_4_lut (.A(new_sboxw[0]), .B(n33506), .C(update_type[0]), 
         .D(n4_adj_7932), .Z(n2_adj_7933)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_64_i2_4_lut.init = 16'h3aca;
    LUT4 mux_626_Mux_69_i2_4_lut (.A(new_sboxw[5]), .B(n7_adj_7934), .C(update_type[0]), 
         .D(n8_adj_7829), .Z(n2_adj_7935)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_69_i2_4_lut.init = 16'h3aca;
    LUT4 mux_626_Mux_76_i2_4_lut (.A(new_sboxw[12]), .B(n5_adj_7936), .C(update_type[0]), 
         .D(n6_adj_7937), .Z(n2_adj_7938)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_76_i2_4_lut.init = 16'h3aca;
    LUT4 mux_626_Mux_84_i2_4_lut (.A(new_sboxw[20]), .B(n5_adj_7907), .C(update_type[0]), 
         .D(n6_adj_7939), .Z(n2_adj_7940)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_84_i2_4_lut.init = 16'h3aca;
    LUT4 i27785_3_lut_4_lut (.A(\block_new_127__N_1645[75] ), .B(update_type[0]), 
         .C(n33844), .D(n13071), .Z(n4540[11])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27785_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_626_Mux_92_i2_4_lut (.A(new_sboxw[28]), .B(n5_adj_7926), .C(update_type[0]), 
         .D(n6_adj_7941), .Z(n2_adj_7942)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_92_i2_4_lut.init = 16'h3aca;
    LUT4 mux_626_Mux_93_i2_4_lut (.A(new_sboxw[29]), .B(n7_adj_7943), .C(update_type[0]), 
         .D(n8_adj_7944), .Z(n2_adj_7945)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_93_i2_4_lut.init = 16'h3aca;
    LUT4 mux_626_Mux_99_i2_4_lut (.A(new_sboxw[3]), .B(n5_adj_7946), .C(update_type[0]), 
         .D(n6_adj_7947), .Z(n2_adj_7948)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_99_i2_4_lut.init = 16'h3aca;
    LUT4 mux_626_Mux_100_i2_4_lut (.A(new_sboxw[4]), .B(n7_adj_7949), .C(update_type[0]), 
         .D(n8_adj_7950), .Z(n2_adj_7951)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_100_i2_4_lut.init = 16'h3aca;
    LUT4 i27587_3_lut_4_lut (.A(block_new_127__N_1645_c[74]), .B(update_type[0]), 
         .C(n33844), .D(n13070), .Z(n4540[10])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27587_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_626_Mux_101_i2_4_lut (.A(new_sboxw[5]), .B(n5_adj_7952), .C(update_type[0]), 
         .D(n6_adj_7953), .Z(n2_adj_7954)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_101_i2_4_lut.init = 16'h3aca;
    LUT4 i2_2_lut_3_lut_4_lut_adj_112 (.A(block_new_127__N_1901[84]), .B(n33704), 
         .C(n33792), .D(n33793), .Z(n7_adj_7943)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i2_2_lut_3_lut_4_lut_adj_112.init = 16'h6996;
    LUT4 mux_626_Mux_108_i2_4_lut (.A(new_sboxw[12]), .B(n5_adj_7955), .C(update_type[0]), 
         .D(n6_adj_7956), .Z(n2_adj_7957)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_108_i2_4_lut.init = 16'h3aca;
    LUT4 i2_2_lut_3_lut_4_lut_adj_113 (.A(block_new_127__N_1901[84]), .B(n33704), 
         .C(n12748), .D(n33793), .Z(n6_adj_7941)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i2_2_lut_3_lut_4_lut_adj_113.init = 16'h6996;
    LUT4 i2_2_lut_3_lut_4_lut_adj_114 (.A(block_new_127__N_1901[110]), .B(block_new_127__N_1901[127]), 
         .C(n33839), .D(block_new_127__N_1901[111]), .Z(n7_adj_7958)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i2_2_lut_3_lut_4_lut_adj_114.init = 16'h6996;
    LUT4 i1_2_lut_rep_275_3_lut_4_lut (.A(block_new_127__N_1901[110]), .B(block_new_127__N_1901[127]), 
         .C(n33756), .D(block_new_127__N_1901[111]), .Z(n33579)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_rep_275_3_lut_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_368_3_lut (.A(block_new_127__N_1901[110]), .B(block_new_127__N_1901[127]), 
         .C(block_new_127__N_1901[111]), .Z(n33672)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_rep_368_3_lut.init = 16'h9696;
    LUT4 block_127__I_0_i122_2_lut (.A(\block_reg[0] [25]), .B(round_key[121]), 
         .Z(\block_new_127__N_1645[121] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i122_2_lut.init = 16'h6666;
    LUT4 i2_2_lut_3_lut_4_lut_adj_115 (.A(block_new_127__N_1901[92]), .B(n33705), 
         .C(n12748), .D(n33792), .Z(n6_adj_7927)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i2_2_lut_3_lut_4_lut_adj_115.init = 16'h6996;
    LUT4 i3_3_lut_4_lut_adj_116 (.A(block_new_127__N_1901[92]), .B(n33705), 
         .C(block_new_127__N_1901[77]), .D(n33804), .Z(n8_adj_7944)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i3_3_lut_4_lut_adj_116.init = 16'h6996;
    LUT4 i27585_3_lut_4_lut (.A(\block_new_127__N_1645[73] ), .B(update_type[0]), 
         .C(n33844), .D(n13069), .Z(n4540[9])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27585_3_lut_4_lut.init = 16'hf808;
    LUT4 i27659_3_lut_4_lut (.A(block_new_127__N_1645_c[72]), .B(update_type[0]), 
         .C(n33844), .D(n13068), .Z(n4540[8])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27659_3_lut_4_lut.init = 16'hf808;
    LUT4 i27231_3_lut_4_lut (.A(block_new_127__N_1645_c[103]), .B(update_type[0]), 
         .C(n33844), .D(n13067), .Z(n4540[7])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27231_3_lut_4_lut.init = 16'hf808;
    LUT4 new_block_127__I_0_i127_2_lut (.A(dec_new_block[126]), .B(round_key[126]), 
         .Z(block_new_127__N_1901[126])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i127_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i112_2_lut (.A(dec_new_block[111]), .B(round_key[111]), 
         .Z(block_new_127__N_1901[111])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i112_2_lut.init = 16'h6666;
    LUT4 i2_2_lut_3_lut_4_lut_adj_117 (.A(n33797), .B(n33705), .C(n33588), 
         .D(n33803), .Z(n6_adj_7953)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i2_2_lut_3_lut_4_lut_adj_117.init = 16'h6996;
    LUT4 i27583_3_lut_4_lut (.A(\block_new_127__N_1645[102] ), .B(update_type[0]), 
         .C(n33844), .D(n13066), .Z(n4540[6])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27583_3_lut_4_lut.init = 16'hf808;
    LUT4 i27735_3_lut_4_lut (.A(block_new_127__N_1645_c[101]), .B(update_type[0]), 
         .C(n33844), .D(n13065), .Z(n4540[5])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27735_3_lut_4_lut.init = 16'hf808;
    LUT4 i2_2_lut_3_lut_4_lut_adj_118 (.A(n33797), .B(n33705), .C(n33702), 
         .D(n33803), .Z(n6_adj_7929)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i2_2_lut_3_lut_4_lut_adj_118.init = 16'h6996;
    LUT4 i27657_3_lut_4_lut (.A(block_new_127__N_1645_c[100]), .B(update_type[0]), 
         .C(n33844), .D(n13064), .Z(n4540[4])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27657_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_626_Mux_5_i2_4_lut (.A(new_sboxw[5]), .B(n33525), .C(update_type[0]), 
         .D(n4_adj_7959), .Z(n2_adj_7960)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_5_i2_4_lut.init = 16'h3aca;
    LUT4 mux_626_Mux_43_i2_4_lut (.A(new_sboxw[11]), .B(n33509), .C(update_type[0]), 
         .D(n4_adj_7961), .Z(n2_adj_7962)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_43_i2_4_lut.init = 16'h3aca;
    LUT4 mux_626_Mux_49_i2_4_lut (.A(new_sboxw[17]), .B(n7_adj_7871), .C(update_type[0]), 
         .D(n8_adj_7963), .Z(n2_adj_7964)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_49_i2_4_lut.init = 16'h3aca;
    LUT4 mux_626_Mux_59_i2_4_lut (.A(new_sboxw[27]), .B(n5_adj_7965), .C(update_type[0]), 
         .D(n6_adj_7966), .Z(n2_adj_7967)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_59_i2_4_lut.init = 16'h3aca;
    LUT4 i1_2_lut_3_lut_adj_119 (.A(block_new_127__N_1901[30]), .B(block_new_127__N_1901[15]), 
         .C(block_new_127__N_1901[23]), .Z(n5_adj_7713)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_3_lut_adj_119.init = 16'h9696;
    LUT4 i1_2_lut_3_lut_adj_120 (.A(block_new_127__N_1901[30]), .B(block_new_127__N_1901[15]), 
         .C(block_new_127__N_1901[7]), .Z(n5_adj_7809)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_3_lut_adj_120.init = 16'h9696;
    LUT4 mux_626_Mux_85_i2_4_lut (.A(new_sboxw[21]), .B(n7_adj_7968), .C(update_type[0]), 
         .D(n8_adj_7969), .Z(n2_adj_7970)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_85_i2_4_lut.init = 16'h3aca;
    LUT4 mux_626_Mux_91_i2_4_lut (.A(new_sboxw[27]), .B(n33507), .C(update_type[0]), 
         .D(n4_adj_7971), .Z(n2_adj_7972)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_91_i2_4_lut.init = 16'h3aca;
    LUT4 mux_626_Mux_105_i2_4_lut (.A(new_sboxw[9]), .B(n7_adj_7973), .C(update_type[0]), 
         .D(n8_adj_7676), .Z(n2_adj_7974)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_105_i2_4_lut.init = 16'h3aca;
    LUT4 mux_626_Mux_107_i2_4_lut (.A(new_sboxw[11]), .B(n7_adj_7975), .C(update_type[0]), 
         .D(n8_adj_7976), .Z(n2_adj_7977)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_107_i2_4_lut.init = 16'h3aca;
    LUT4 i3_3_lut_4_lut_adj_121 (.A(block_new_127__N_1901[125]), .B(n33710), 
         .C(block_new_127__N_1901[118]), .D(n29339), .Z(n8_adj_7789)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i3_3_lut_4_lut_adj_121.init = 16'h6996;
    LUT4 mux_626_Mux_115_i2_4_lut (.A(new_sboxw[19]), .B(n5_adj_7978), .C(update_type[0]), 
         .D(n6_adj_7979), .Z(n2_adj_7980)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_115_i2_4_lut.init = 16'h3aca;
    LUT4 new_block_127__I_0_i122_2_lut (.A(dec_new_block[121]), .B(round_key[121]), 
         .Z(block_new_127__N_1901[121])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i122_2_lut.init = 16'h6666;
    LUT4 i27655_3_lut_4_lut (.A(\block_new_127__N_1645[99] ), .B(update_type[0]), 
         .C(n33844), .D(n13063), .Z(n4540[3])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27655_3_lut_4_lut.init = 16'hf808;
    LUT4 i27581_3_lut_4_lut (.A(\block_new_127__N_1645[98] ), .B(update_type[0]), 
         .C(n33844), .D(n13062), .Z(n4540[2])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27581_3_lut_4_lut.init = 16'hf808;
    LUT4 i1_2_lut_4_lut_adj_122 (.A(block_new_127__N_1901[79]), .B(n33708), 
         .C(block_new_127__N_1901[94]), .D(block_new_127__N_1901[86]), .Z(n4_adj_7858)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_4_lut_adj_122.init = 16'h6996;
    LUT4 i3_3_lut_4_lut_adj_123 (.A(block_new_127__N_1901[101]), .B(n33710), 
         .C(block_new_127__N_1901[116]), .D(block_new_127__N_1901[125]), 
         .Z(n8_adj_7969)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i3_3_lut_4_lut_adj_123.init = 16'h6996;
    LUT4 i1_2_lut_3_lut_adj_124 (.A(block_new_127__N_1901[121]), .B(block_new_127__N_1901[96]), 
         .C(n33791), .Z(n5_adj_7695)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_3_lut_adj_124.init = 16'h9696;
    LUT4 i27507_3_lut_4_lut (.A(\block_new_127__N_1645[97] ), .B(update_type[0]), 
         .C(n33844), .D(n13061), .Z(n4540[1])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27507_3_lut_4_lut.init = 16'hf808;
    LUT4 i3_3_lut_4_lut_adj_125 (.A(block_new_127__N_1901[98]), .B(block_new_127__N_1901[122]), 
         .C(block_new_127__N_1901[114]), .D(n33767), .Z(n8_adj_7824)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i3_3_lut_4_lut_adj_125.init = 16'h6996;
    PFUMX i9324 (.BLUT(n14933), .ALUT(n14934), .C0(n30080), .Z(round_ctr_new_c[2]));
    LUT4 i2_3_lut_rep_372_4_lut (.A(block_new_127__N_1901[47]), .B(block_new_127__N_1901[46]), 
         .C(block_new_127__N_1901[54]), .D(block_new_127__N_1901[63]), .Z(n33676)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i2_3_lut_rep_372_4_lut.init = 16'h6996;
    LUT4 i3_2_lut_3_lut (.A(block_new_127__N_1901[38]), .B(block_new_127__N_1901[62]), 
         .C(n29390), .Z(n9_adj_7830)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i3_2_lut_3_lut.init = 16'h9696;
    LUT4 i2_2_lut_3_lut_4_lut_adj_126 (.A(block_new_127__N_1901[38]), .B(block_new_127__N_1901[62]), 
         .C(n33684), .D(n33800), .Z(n6_adj_7743)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i2_2_lut_3_lut_4_lut_adj_126.init = 16'h6996;
    LUT4 i2_3_lut_rep_373_4_lut (.A(block_new_127__N_1901[5]), .B(block_new_127__N_1901[4]), 
         .C(block_new_127__N_1901[12]), .D(block_new_127__N_1901[21]), .Z(n33677)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i2_3_lut_rep_373_4_lut.init = 16'h6996;
    LUT4 i3_2_lut_3_lut_adj_127 (.A(block_new_127__N_1901[5]), .B(block_new_127__N_1901[4]), 
         .C(n29143), .Z(n9_adj_7817)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i3_2_lut_3_lut_adj_127.init = 16'h9696;
    LUT4 i1_2_lut_3_lut_4_lut_adj_128 (.A(block_new_127__N_1901[70]), .B(block_new_127__N_1901[94]), 
         .C(block_new_127__N_1901[89]), .D(block_new_127__N_1901[74]), .Z(n5_adj_7853)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_3_lut_4_lut_adj_128.init = 16'h6996;
    LUT4 i2_2_lut_rep_378_3_lut (.A(block_new_127__N_1901[70]), .B(block_new_127__N_1901[94]), 
         .C(block_new_127__N_1901[74]), .Z(n33682)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i2_2_lut_rep_378_3_lut.init = 16'h9696;
    LUT4 i2_2_lut_3_lut (.A(block_new_127__N_1901[70]), .B(block_new_127__N_1901[94]), 
         .C(block_new_127__N_1901[90]), .Z(n7_adj_7794)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i2_2_lut_3_lut.init = 16'h9696;
    LUT4 i1_2_lut_3_lut_adj_129 (.A(block_new_127__N_1901[70]), .B(block_new_127__N_1901[94]), 
         .C(block_new_127__N_1901[87]), .Z(n5_adj_7769)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_3_lut_adj_129.init = 16'h9696;
    LUT4 i2_2_lut_3_lut_4_lut_adj_130 (.A(block_new_127__N_1901[69]), .B(block_new_127__N_1901[94]), 
         .C(n33793), .D(n33792), .Z(n6_adj_7797)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i2_2_lut_3_lut_4_lut_adj_130.init = 16'h6996;
    LUT4 i1_2_lut_rep_365_3_lut_4_lut (.A(block_new_127__N_1901[86]), .B(block_new_127__N_1901[78]), 
         .C(block_new_127__N_1901[95]), .D(block_new_127__N_1901[79]), .Z(n33669)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_365_3_lut_4_lut.init = 16'h6996;
    LUT4 i2_2_lut_3_lut_4_lut_adj_131 (.A(block_new_127__N_1901[86]), .B(block_new_127__N_1901[78]), 
         .C(block_new_127__N_1901[94]), .D(block_new_127__N_1901[69]), .Z(n7_adj_7860)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i2_2_lut_3_lut_4_lut_adj_131.init = 16'h6996;
    LUT4 i3_2_lut_3_lut_4_lut_adj_132 (.A(block_new_127__N_1901[21]), .B(n33784), 
         .C(n33828), .D(n33686), .Z(n9_adj_7707)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i3_2_lut_3_lut_4_lut_adj_132.init = 16'h6996;
    LUT4 i2_3_lut_rep_380_4_lut (.A(block_new_127__N_1901[44]), .B(block_new_127__N_1901[36]), 
         .C(block_new_127__N_1901[37]), .D(block_new_127__N_1901[53]), .Z(n33684)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i2_3_lut_rep_380_4_lut.init = 16'h6996;
    LUT4 i1_4_lut_adj_133 (.A(dec_ctrl_new_2__N_2032), .B(n33842), .C(n20699), 
         .D(n33844), .Z(block_w3_we)) /* synthesis lut_function=(!(A+!(B (C+(D))+!B !((D)+!C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(462[7] 518[14])
    defparam i1_4_lut_adj_133.init = 16'h4450;
    LUT4 i2_3_lut_4_lut (.A(block_new_127__N_1901[46]), .B(block_new_127__N_1901[55]), 
         .C(block_new_127__N_1901[50]), .D(block_new_127__N_1901[56]), .Z(n29393)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i2_3_lut_4_lut.init = 16'h6996;
    LUT4 i2_2_lut_3_lut_4_lut_adj_134 (.A(block_new_127__N_1901[21]), .B(n33784), 
         .C(n33826), .D(n33686), .Z(n6_adj_7778)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i2_2_lut_3_lut_4_lut_adj_134.init = 16'h6996;
    LUT4 i1_2_lut_3_lut_adj_135 (.A(block_new_127__N_1901[46]), .B(block_new_127__N_1901[55]), 
         .C(block_new_127__N_1901[38]), .Z(n5_adj_7864)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_3_lut_adj_135.init = 16'h9696;
    LUT4 i3_2_lut_3_lut_adj_136 (.A(block_new_127__N_1901[14]), .B(block_new_127__N_1901[7]), 
         .C(block_new_127__N_1901[16]), .Z(n9_adj_7866)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i3_2_lut_3_lut_adj_136.init = 16'h9696;
    LUT4 i1_2_lut_3_lut_adj_137 (.A(block_new_127__N_1901[14]), .B(block_new_127__N_1901[7]), 
         .C(block_new_127__N_1901[24]), .Z(n5_adj_7981)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_3_lut_adj_137.init = 16'h9696;
    LUT4 i1_2_lut_3_lut_4_lut_adj_138 (.A(block_new_127__N_1901[14]), .B(block_new_127__N_1901[7]), 
         .C(block_new_127__N_1901[6]), .D(block_new_127__N_1901[31]), .Z(n4_adj_7748)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_3_lut_4_lut_adj_138.init = 16'h6996;
    LUT4 block_127__I_0_i121_2_lut (.A(\block_reg[0] [24]), .B(round_key[120]), 
         .Z(block_new_127__N_1645_c[120])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i121_2_lut.init = 16'h6666;
    LUT4 mux_626_Mux_11_i2_4_lut (.A(new_sboxw[11]), .B(n5_adj_7982), .C(update_type[0]), 
         .D(n6), .Z(n2_adj_7983)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_11_i2_4_lut.init = 16'h3aca;
    LUT4 mux_626_Mux_27_i2_4_lut (.A(new_sboxw[27]), .B(n7_adj_7984), .C(update_type[0]), 
         .D(n8_adj_7985), .Z(n2_adj_7986)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_27_i2_4_lut.init = 16'h3aca;
    LUT4 mux_626_Mux_51_i2_4_lut (.A(new_sboxw[19]), .B(n9_adj_7987), .C(update_type[0]), 
         .D(n10_adj_7988), .Z(n2_adj_7989)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_51_i2_4_lut.init = 16'h3aca;
    LUT4 i1_2_lut_3_lut_adj_139 (.A(block_new_127__N_1901[9]), .B(block_new_127__N_1901[1]), 
         .C(block_new_127__N_1901[26]), .Z(n4_adj_7839)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_3_lut_adj_139.init = 16'h9696;
    LUT4 i1_2_lut_4_lut_adj_140 (.A(block_new_127__N_1901[4]), .B(n33780), 
         .C(block_new_127__N_1901[28]), .D(block_new_127__N_1901[21]), .Z(n4_adj_7814)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_4_lut_adj_140.init = 16'h6996;
    LUT4 i1_2_lut_3_lut_4_lut_adj_141 (.A(block_new_127__N_1901[102]), .B(block_new_127__N_1901[118]), 
         .C(n33767), .D(n33791), .Z(n4_adj_7750)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_3_lut_4_lut_adj_141.init = 16'h6996;
    LUT4 i1_2_lut_rep_279_3_lut_4_lut (.A(block_new_127__N_1901[102]), .B(block_new_127__N_1901[118]), 
         .C(block_new_127__N_1901[106]), .D(block_new_127__N_1901[126]), 
         .Z(n33583)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_279_3_lut_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_384_3_lut (.A(block_new_127__N_1901[102]), .B(block_new_127__N_1901[118]), 
         .C(block_new_127__N_1901[126]), .Z(n33688)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_384_3_lut.init = 16'h9696;
    LUT4 mux_626_Mux_75_i2_4_lut (.A(new_sboxw[11]), .B(n5_adj_7990), .C(update_type[0]), 
         .D(n6_adj_7768), .Z(n2_adj_7991)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_75_i2_4_lut.init = 16'h3aca;
    LUT4 mux_626_Mux_83_i2_4_lut (.A(new_sboxw[19]), .B(n7_adj_7992), .C(update_type[0]), 
         .D(n8_adj_7674), .Z(n2_adj_7993)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_83_i2_4_lut.init = 16'h3aca;
    LUT4 mux_626_Mux_123_i2_4_lut (.A(new_sboxw[27]), .B(n5_adj_7994), .C(update_type[0]), 
         .D(n6_adj_7816), .Z(n2_adj_7995)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_123_i2_4_lut.init = 16'h3aca;
    LUT4 i2_2_lut_3_lut_4_lut_adj_142 (.A(block_new_127__N_1901[102]), .B(block_new_127__N_1901[118]), 
         .C(n33830), .D(n33791), .Z(n7_adj_7782)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i2_2_lut_3_lut_4_lut_adj_142.init = 16'h6996;
    LUT4 mux_626_Mux_125_i2_4_lut (.A(new_sboxw[29]), .B(n7_adj_7996), .C(update_type[0]), 
         .D(n8_adj_7688), .Z(n2_adj_7997)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_125_i2_4_lut.init = 16'h3aca;
    LUT4 new_block_127__I_0_i121_2_lut (.A(dec_new_block[120]), .B(round_key[120]), 
         .Z(block_new_127__N_1901[120])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i121_2_lut.init = 16'h6666;
    LUT4 i1_4_lut_rep_542 (.A(n6347[3]), .B(n6347[1]), .C(n6347[2]), .D(n33848), 
         .Z(n33846)) /* synthesis lut_function=(!(A+!(B (C)+!B (C+!(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_encipher_block.v(164[17:30])
    defparam i1_4_lut_rep_542.init = 16'h5051;
    LUT4 i1_2_lut_rep_385_3_lut (.A(block_new_127__N_1901[119]), .B(block_new_127__N_1901[120]), 
         .C(block_new_127__N_1901[113]), .Z(n33689)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_385_3_lut.init = 16'h9696;
    LUT4 i14475_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[3]), .Z(n13063)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14475_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i15180_3_lut_4_lut (.A(n33849), .B(n33935), .C(n6362[2]), .D(update_type[0]), 
         .Z(n20702)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (D)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i15180_3_lut_4_lut.init = 16'hff20;
    LUT4 i14474_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[4]), .Z(n13064)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14474_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14473_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[5]), .Z(n13065)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14473_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14472_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[6]), .Z(n13066)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14472_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14471_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[7]), .Z(n13067)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14471_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i15177_3_lut_4_lut (.A(n33849), .B(n33935), .C(n6362[3]), .D(update_type[0]), 
         .Z(n20699)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (D)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i15177_3_lut_4_lut.init = 16'hff20;
    LUT4 i14477_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[1]), .Z(n13061)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14477_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i1_2_lut_rep_374_3_lut (.A(block_new_127__N_1901[103]), .B(block_new_127__N_1901[104]), 
         .C(block_new_127__N_1901[97]), .Z(n33678)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_rep_374_3_lut.init = 16'h9696;
    LUT4 i14470_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[8]), .Z(n13068)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14470_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14469_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[9]), .Z(n13069)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14469_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14468_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[10]), .Z(n13070)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14468_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14467_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[11]), .Z(n13071)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14467_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14466_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[12]), .Z(n13072)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14466_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14465_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[13]), .Z(n13073)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14465_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14464_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[14]), .Z(n13074)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14464_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14463_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[15]), .Z(n13075)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14463_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i1_2_lut_3_lut_4_lut_adj_143 (.A(block_new_127__N_1901[103]), .B(block_new_127__N_1901[104]), 
         .C(block_new_127__N_1901[113]), .D(block_new_127__N_1901[97]), 
         .Z(n5_adj_7821)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_3_lut_4_lut_adj_143.init = 16'h6996;
    LUT4 i15186_3_lut_4_lut (.A(n33849), .B(n33935), .C(n6362[0]), .D(update_type[0]), 
         .Z(n20708)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (D)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i15186_3_lut_4_lut.init = 16'hff20;
    LUT4 i14462_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[16]), .Z(n13076)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14462_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14461_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[17]), .Z(n13077)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14461_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14460_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[18]), .Z(n13078)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14460_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14459_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[19]), .Z(n13079)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14459_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i15183_3_lut_4_lut (.A(n33849), .B(n33935), .C(n6362[1]), .D(update_type[0]), 
         .Z(n20705)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (D)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i15183_3_lut_4_lut.init = 16'hff20;
    LUT4 i14458_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[20]), .Z(n13080)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14458_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14457_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[21]), .Z(n13081)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14457_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14456_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[22]), .Z(n13082)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14456_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14455_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[23]), .Z(n13083)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14455_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i1_2_lut_4_lut_adj_144 (.A(n33760), .B(block_new_127__N_1901[63]), 
         .C(block_new_127__N_1901[54]), .D(block_new_127__N_1901[39]), .Z(n4_adj_7998)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_4_lut_adj_144.init = 16'h6996;
    LUT4 i14454_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[24]), .Z(n13084)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14454_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14453_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[25]), .Z(n13085)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14453_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14452_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[26]), .Z(n13086)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14452_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14451_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[27]), .Z(n13087)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14451_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14450_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[28]), .Z(n13088)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14450_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14449_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[29]), .Z(n13089)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14449_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14448_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[30]), .Z(n13090)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14448_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14447_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[31]), .Z(n13091)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14447_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14446_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[32]), .Z(n13092)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14446_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14445_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[33]), .Z(n13093)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14445_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14444_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[34]), .Z(n13094)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14444_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14443_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[35]), .Z(n13095)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14443_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i2_2_lut_3_lut_4_lut_adj_145 (.A(block_new_127__N_1901[109]), .B(block_new_127__N_1901[108]), 
         .C(n33714), .D(n33839), .Z(n7_adj_7880)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i2_2_lut_3_lut_4_lut_adj_145.init = 16'h6996;
    LUT4 i14442_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[36]), .Z(n13096)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14442_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14441_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[37]), .Z(n13097)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14441_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14440_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[38]), .Z(n13098)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14440_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14439_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[39]), .Z(n13099)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14439_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i1_2_lut_rep_387_3_lut (.A(block_new_127__N_1901[109]), .B(block_new_127__N_1901[108]), 
         .C(block_new_127__N_1901[124]), .Z(n33691)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_rep_387_3_lut.init = 16'h9696;
    LUT4 i14438_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[40]), .Z(n13100)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14438_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14437_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[41]), .Z(n13101)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14437_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14436_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[42]), .Z(n13102)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14436_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14435_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[43]), .Z(n13103)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14435_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i1_2_lut_3_lut_adj_146 (.A(block_new_127__N_1901[64]), .B(block_new_127__N_1901[80]), 
         .C(block_new_127__N_1901[88]), .Z(n4_adj_7893)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_3_lut_adj_146.init = 16'h9696;
    LUT4 i14434_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[44]), .Z(n13104)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14434_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14433_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[45]), .Z(n13105)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14433_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14432_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[46]), .Z(n13106)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14432_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14431_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[47]), .Z(n13107)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14431_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14430_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[48]), .Z(n13108)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14430_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14429_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[49]), .Z(n13109)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14429_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14428_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[50]), .Z(n13110)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14428_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14427_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[51]), .Z(n13111)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14427_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14426_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[52]), .Z(n13112)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14426_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14425_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[53]), .Z(n13113)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14425_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14424_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[54]), .Z(n13114)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14424_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14423_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[55]), .Z(n13115)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14423_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14422_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[56]), .Z(n13116)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14422_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14421_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[57]), .Z(n13117)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14421_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14420_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[58]), .Z(n13118)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14420_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i1_2_lut_rep_389_3_lut (.A(block_new_127__N_1901[47]), .B(block_new_127__N_1901[56]), 
         .C(block_new_127__N_1901[55]), .Z(n33693)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_389_3_lut.init = 16'h9696;
    LUT4 i2_2_lut_3_lut_4_lut_adj_147 (.A(block_new_127__N_1901[47]), .B(block_new_127__N_1901[56]), 
         .C(block_new_127__N_1901[49]), .D(block_new_127__N_1901[55]), .Z(n7_adj_7732)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i2_2_lut_3_lut_4_lut_adj_147.init = 16'h6996;
    LUT4 i14419_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[59]), .Z(n13119)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14419_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14418_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[60]), .Z(n13120)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14418_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14417_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[61]), .Z(n13121)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14417_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14416_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[62]), .Z(n13122)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14416_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14415_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[63]), .Z(n13123)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14415_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14414_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[64]), .Z(n13124)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14414_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14413_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[65]), .Z(n13125)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14413_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14412_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[66]), .Z(n13126)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14412_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i1_2_lut_rep_391_3_lut (.A(block_new_127__N_1901[14]), .B(block_new_127__N_1901[22]), 
         .C(block_new_127__N_1901[7]), .Z(n33695)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_391_3_lut.init = 16'h9696;
    LUT4 i14411_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[67]), .Z(n13127)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14411_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14410_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[68]), .Z(n13128)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14410_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14409_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[69]), .Z(n13129)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14409_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14408_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[70]), .Z(n13130)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14408_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i2_3_lut_rep_364_4_lut (.A(block_new_127__N_1901[14]), .B(block_new_127__N_1901[22]), 
         .C(block_new_127__N_1901[26]), .D(block_new_127__N_1901[10]), .Z(n33668)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i2_3_lut_rep_364_4_lut.init = 16'h6996;
    LUT4 i14407_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[71]), .Z(n13131)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14407_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14406_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[72]), .Z(n13132)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14406_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14405_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[73]), .Z(n13133)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14405_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14404_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[74]), .Z(n13134)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14404_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i1_2_lut_3_lut_adj_148 (.A(block_new_127__N_1901[23]), .B(block_new_127__N_1901[24]), 
         .C(block_new_127__N_1901[0]), .Z(n5_adj_7777)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_3_lut_adj_148.init = 16'h9696;
    LUT4 i2_3_lut_rep_472 (.A(block_new_127__N_1901[18]), .B(block_new_127__N_1901[6]), 
         .C(block_new_127__N_1901[30]), .Z(n33776)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i2_3_lut_rep_472.init = 16'h9696;
    LUT4 i14403_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[75]), .Z(n13135)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14403_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i1_2_lut_4_lut_adj_149 (.A(block_new_127__N_1901[18]), .B(block_new_127__N_1901[6]), 
         .C(block_new_127__N_1901[30]), .D(block_new_127__N_1901[8]), .Z(n6_adj_7999)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_4_lut_adj_149.init = 16'h6996;
    LUT4 i14402_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[76]), .Z(n13136)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14402_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14401_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[77]), .Z(n13137)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14401_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14400_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[78]), .Z(n13138)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14400_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14399_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[79]), .Z(n13139)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14399_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i2_2_lut_3_lut_4_lut_adj_150 (.A(block_new_127__N_1901[44]), .B(n33799), 
         .C(n33706), .D(n33699), .Z(n6_adj_7804)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i2_2_lut_3_lut_4_lut_adj_150.init = 16'h6996;
    LUT4 i14398_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[80]), .Z(n13140)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14398_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14397_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[81]), .Z(n13141)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14397_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14396_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[82]), .Z(n13142)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14396_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14395_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[83]), .Z(n13143)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14395_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14394_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[84]), .Z(n13144)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14394_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14393_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[85]), .Z(n13145)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14393_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14392_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[86]), .Z(n13146)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14392_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i3_2_lut_3_lut_4_lut_adj_151 (.A(block_new_127__N_1901[25]), .B(block_new_127__N_1901[17]), 
         .C(block_new_127__N_1901[8]), .D(block_new_127__N_1901[31]), .Z(n9_adj_7745)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i3_2_lut_3_lut_4_lut_adj_151.init = 16'h6996;
    LUT4 i14391_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[87]), .Z(n13147)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14391_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14390_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[88]), .Z(n13148)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14390_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14389_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[89]), .Z(n13149)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14389_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i1_2_lut_3_lut_adj_152 (.A(block_new_127__N_1901[19]), .B(block_new_127__N_1901[23]), 
         .C(n12810), .Z(n5_adj_7908)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_3_lut_adj_152.init = 16'h9696;
    LUT4 i14388_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[90]), .Z(n13150)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14388_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14387_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[91]), .Z(n13151)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14387_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14386_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[92]), .Z(n13152)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14386_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14385_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[93]), .Z(n13153)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14385_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14384_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[94]), .Z(n13154)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14384_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14383_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[95]), .Z(n13155)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14383_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14382_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[96]), .Z(n13156)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14382_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14381_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[97]), .Z(n13157)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14381_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i1_2_lut_rep_280_3_lut_4_lut (.A(block_new_127__N_1901[5]), .B(block_new_127__N_1901[21]), 
         .C(block_new_127__N_1901[30]), .D(n33780), .Z(n33584)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_rep_280_3_lut_4_lut.init = 16'h6996;
    LUT4 i14380_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[98]), .Z(n13158)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14380_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14379_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[99]), .Z(n13159)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14379_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14378_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[100]), .Z(n13160)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14378_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14377_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[101]), .Z(n13161)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14377_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14376_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[102]), .Z(n13162)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14376_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14375_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[103]), .Z(n13163)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14375_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14374_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[104]), .Z(n13164)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14374_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14373_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[105]), .Z(n13165)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14373_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14372_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[106]), .Z(n13166)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14372_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14371_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[107]), .Z(n13167)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14371_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i2_3_lut_rep_370_4_lut (.A(block_new_127__N_1901[29]), .B(block_new_127__N_1901[13]), 
         .C(block_new_127__N_1901[28]), .D(block_new_127__N_1901[4]), .Z(n33674)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i2_3_lut_rep_370_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_382_3_lut (.A(block_new_127__N_1901[29]), .B(block_new_127__N_1901[13]), 
         .C(block_new_127__N_1901[5]), .Z(n33686)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_382_3_lut.init = 16'h9696;
    LUT4 i14370_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[108]), .Z(n13168)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14370_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14369_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[109]), .Z(n13169)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14369_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14368_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[110]), .Z(n13170)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14368_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14367_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[111]), .Z(n13171)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14367_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14366_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[112]), .Z(n13172)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14366_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i1_2_lut_rep_535_4_lut (.A(dec_new_block[100]), .B(round_key[100]), 
         .C(dec_new_block[116]), .D(round_key[116]), .Z(n33839)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_rep_535_4_lut.init = 16'h6996;
    LUT4 i14365_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[113]), .Z(n13173)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14365_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14364_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[114]), .Z(n13174)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14364_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14363_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[115]), .Z(n13175)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14363_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i1_2_lut_3_lut_4_lut_adj_153 (.A(block_new_127__N_1901[29]), .B(block_new_127__N_1901[13]), 
         .C(n33782), .D(block_new_127__N_1901[5]), .Z(n4_adj_7872)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_3_lut_4_lut_adj_153.init = 16'h6996;
    LUT4 i14362_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[116]), .Z(n13176)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14362_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14361_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[117]), .Z(n13177)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14361_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14360_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[118]), .Z(n13178)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14360_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14359_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[119]), .Z(n13179)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14359_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14358_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[120]), .Z(n13180)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14358_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i3_3_lut_4_lut_adj_154 (.A(block_new_127__N_1901[17]), .B(block_new_127__N_1901[9]), 
         .C(block_new_127__N_1901[25]), .D(n33825), .Z(n8_adj_7913)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i3_3_lut_4_lut_adj_154.init = 16'h6996;
    LUT4 i14357_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[121]), .Z(n13181)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14357_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14356_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[122]), .Z(n13182)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14356_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14355_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[123]), .Z(n13183)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14355_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14354_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[124]), .Z(n13184)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14354_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i15417_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[0]), .Z(n12933)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i15417_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14351_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[127]), .Z(n13187)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14351_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i2_2_lut_3_lut_4_lut_adj_155 (.A(block_new_127__N_1901[20]), .B(block_new_127__N_1901[12]), 
         .C(n29291), .D(n33783), .Z(n6_adj_7909)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i2_2_lut_3_lut_4_lut_adj_155.init = 16'h6996;
    LUT4 i14476_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[2]), .Z(n13062)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14476_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i14353_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[125]), .Z(n13185)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14353_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i2_2_lut_3_lut_4_lut_adj_156 (.A(block_new_127__N_1901[20]), .B(block_new_127__N_1901[12]), 
         .C(n29288), .D(n33783), .Z(n6_adj_7919)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i2_2_lut_3_lut_4_lut_adj_156.init = 16'h6996;
    LUT4 i14352_2_lut_3_lut_3_lut_4_lut (.A(n33849), .B(n33935), .C(update_type[0]), 
         .D(block_new_127__N_1901[126]), .Z(n13186)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i14352_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i2_2_lut_3_lut_4_lut_adj_157 (.A(block_new_127__N_1901[44]), .B(n33799), 
         .C(n33699), .D(n4770[4]), .Z(n6_adj_7837)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i2_2_lut_3_lut_4_lut_adj_157.init = 16'h6996;
    LUT4 i2_3_lut_rep_278_4_lut (.A(block_new_127__N_1901[39]), .B(n33812), 
         .C(n33800), .D(n33763), .Z(n33582)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i2_3_lut_rep_278_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_285_3_lut_4_lut (.A(block_new_127__N_1901[99]), .B(block_new_127__N_1901[103]), 
         .C(block_new_127__N_1901[125]), .D(n33808), .Z(n33589)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_285_3_lut_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_406_3_lut_4_lut (.A(block_new_127__N_1901[115]), .B(block_new_127__N_1901[119]), 
         .C(block_new_127__N_1901[103]), .D(block_new_127__N_1901[99]), 
         .Z(n33710)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_406_3_lut_4_lut.init = 16'h6996;
    LUT4 block_127__I_0_i71_2_lut (.A(\block_reg[1] [6]), .B(round_key[70]), 
         .Z(\block_new_127__N_1645[70] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i71_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i70_2_lut (.A(\block_reg[1] [5]), .B(round_key[69]), 
         .Z(\block_new_127__N_1645[69] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i70_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i69_2_lut (.A(\block_reg[1] [4]), .B(round_key[68]), 
         .Z(\block_new_127__N_1645[68] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i69_2_lut.init = 16'h6666;
    LUT4 i3_3_lut_4_lut_adj_158 (.A(block_new_127__N_1901[115]), .B(block_new_127__N_1901[119]), 
         .C(n33837), .D(n29444), .Z(n8_adj_7881)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i3_3_lut_4_lut_adj_158.init = 16'h6996;
    LUT4 i3_2_lut_3_lut_4_lut_adj_159 (.A(block_new_127__N_1901[44]), .B(n33799), 
         .C(n33700), .D(n33798), .Z(n9_adj_7735)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i3_2_lut_3_lut_4_lut_adj_159.init = 16'h6996;
    LUT4 i2_3_lut_rep_276_4_lut (.A(block_new_127__N_1901[20]), .B(block_new_127__N_1901[12]), 
         .C(block_new_127__N_1901[23]), .D(n33674), .Z(n33580)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i2_3_lut_rep_276_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_3_lut_4_lut_adj_160 (.A(block_new_127__N_1901[27]), .B(block_new_127__N_1901[31]), 
         .C(n33677), .D(block_new_127__N_1901[29]), .Z(n4_adj_7841)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_3_lut_4_lut_adj_160.init = 16'h6996;
    LUT4 i1_2_lut_rep_383_3_lut (.A(block_new_127__N_1901[27]), .B(block_new_127__N_1901[31]), 
         .C(block_new_127__N_1901[30]), .Z(n33687)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_383_3_lut.init = 16'h9696;
    LUT4 i2_2_lut_3_lut_adj_161 (.A(block_new_127__N_1901[27]), .B(block_new_127__N_1901[31]), 
         .C(block_new_127__N_1901[13]), .Z(n7_adj_7911)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i2_2_lut_3_lut_adj_161.init = 16'h9696;
    LUT4 i2_2_lut_3_lut_4_lut_adj_162 (.A(block_new_127__N_1901[29]), .B(n33783), 
         .C(n11918), .D(n33788), .Z(n6_adj_7807)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i2_2_lut_3_lut_4_lut_adj_162.init = 16'h6996;
    LUT4 i1_2_lut_3_lut_4_lut_adj_163 (.A(block_new_127__N_1901[27]), .B(block_new_127__N_1901[31]), 
         .C(n33784), .D(block_new_127__N_1901[30]), .Z(n5_adj_7844)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_3_lut_4_lut_adj_163.init = 16'h6996;
    LUT4 i2_3_lut_rep_393_4_lut (.A(block_new_127__N_1901[22]), .B(block_new_127__N_1901[6]), 
         .C(n33823), .D(n33817), .Z(n33697)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i2_3_lut_rep_393_4_lut.init = 16'h6996;
    LUT4 block_127__I_0_i24_2_lut (.A(\block_reg[3] [23]), .B(round_key[23]), 
         .Z(block_new_127__N_1645_c[23])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i24_2_lut.init = 16'h6666;
    LUT4 i1_2_lut_rep_270_4_lut (.A(n33761), .B(block_new_127__N_1901[21]), 
         .C(block_new_127__N_1901[12]), .D(n12090), .Z(n33574)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_rep_270_4_lut.init = 16'h6996;
    LUT4 i27850_2_lut_rep_538_2_lut_3_lut_4_lut (.A(n6363[1]), .B(n33856), 
         .C(update_type[0]), .D(n33935), .Z(n33842)) /* synthesis lut_function=(!(A (C+!(D))+!A (B (C+!(D))+!B (C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i27850_2_lut_rep_538_2_lut_3_lut_4_lut.init = 16'h0f01;
    LUT4 i1_2_lut_rep_369_3_lut (.A(block_new_127__N_1901[22]), .B(block_new_127__N_1901[6]), 
         .C(block_new_127__N_1901[21]), .Z(n33673)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_rep_369_3_lut.init = 16'h9696;
    LUT4 i2_3_lut_4_lut_4_lut_3_lut_4_lut (.A(n6363[1]), .B(n33856), .C(n33935), 
         .D(update_type[0]), .Z(n25333)) /* synthesis lut_function=(A (C+(D))+!A ((C+(D))+!B)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i2_3_lut_4_lut_4_lut_3_lut_4_lut.init = 16'hfff1;
    LUT4 i1_2_lut_3_lut_4_lut_adj_164 (.A(block_new_127__N_1901[22]), .B(block_new_127__N_1901[6]), 
         .C(block_new_127__N_1901[14]), .D(block_new_127__N_1901[21]), .Z(n5_adj_7806)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_3_lut_4_lut_adj_164.init = 16'h6996;
    LUT4 i1_2_lut_3_lut_4_lut_adj_165 (.A(block_new_127__N_1901[76]), .B(block_new_127__N_1901[68]), 
         .C(n33704), .D(n33804), .Z(n5_adj_7696)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_3_lut_4_lut_adj_165.init = 16'h6996;
    LUT4 i1_2_lut_rep_274_3_lut_4_lut (.A(block_new_127__N_1901[76]), .B(block_new_127__N_1901[68]), 
         .C(n33794), .D(n33804), .Z(n33578)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_rep_274_3_lut_4_lut.init = 16'h6996;
    LUT4 i2_3_lut_4_lut_adj_166 (.A(block_new_127__N_1901[76]), .B(block_new_127__N_1901[68]), 
         .C(block_new_127__N_1901[87]), .D(n33794), .Z(n29244)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i2_3_lut_4_lut_adj_166.init = 16'h6996;
    LUT4 i3_3_lut_rep_395_4_lut (.A(block_new_127__N_1901[38]), .B(block_new_127__N_1901[54]), 
         .C(n33806), .D(n5085[3]), .Z(n33699)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i3_3_lut_rep_395_4_lut.init = 16'h6996;
    LUT4 i3_3_lut_4_lut_adj_167 (.A(block_new_127__N_1901[38]), .B(block_new_127__N_1901[54]), 
         .C(block_new_127__N_1901[41]), .D(n33575), .Z(n8_adj_7733)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i3_3_lut_4_lut_adj_167.init = 16'h6996;
    LUT4 i1_2_lut_rep_367_3_lut (.A(block_new_127__N_1901[38]), .B(block_new_127__N_1901[54]), 
         .C(block_new_127__N_1901[62]), .Z(n33671)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_367_3_lut.init = 16'h9696;
    LUT4 i1_2_lut_rep_396_3_lut (.A(block_new_127__N_1901[51]), .B(block_new_127__N_1901[55]), 
         .C(block_new_127__N_1901[60]), .Z(n33700)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_396_3_lut.init = 16'h9696;
    LUT4 i2_2_lut_3_lut_4_lut_adj_168 (.A(block_new_127__N_1901[51]), .B(block_new_127__N_1901[55]), 
         .C(block_new_127__N_1901[36]), .D(block_new_127__N_1901[60]), .Z(n7_adj_7934)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i2_2_lut_3_lut_4_lut_adj_168.init = 16'h6996;
    LUT4 i1_2_lut_rep_371_3_lut (.A(block_new_127__N_1901[51]), .B(block_new_127__N_1901[55]), 
         .C(block_new_127__N_1901[52]), .Z(n33675)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_371_3_lut.init = 16'h9696;
    LUT4 i2_3_lut_4_lut_adj_169 (.A(block_new_127__N_1901[13]), .B(block_new_127__N_1901[5]), 
         .C(n6228[3]), .D(n6327[3]), .Z(n8_adj_8000)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i2_3_lut_4_lut_adj_169.init = 16'h6996;
    LUT4 i2_2_lut_3_lut_4_lut_adj_170 (.A(block_new_127__N_1901[13]), .B(block_new_127__N_1901[5]), 
         .C(n11918), .D(n33788), .Z(n6_adj_7845)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i2_2_lut_3_lut_4_lut_adj_170.init = 16'h6996;
    LUT4 i1_2_lut_rep_215_3_lut_4_lut (.A(block_new_127__N_1901[11]), .B(block_new_127__N_1901[15]), 
         .C(n33697), .D(n12810), .Z(n33519)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_215_3_lut_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_283_3_lut (.A(block_new_127__N_1901[11]), .B(block_new_127__N_1901[15]), 
         .C(n12810), .Z(n33587)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_283_3_lut.init = 16'h9696;
    LUT4 i1_2_lut_3_lut_4_lut_adj_171 (.A(block_new_127__N_1901[11]), .B(block_new_127__N_1901[15]), 
         .C(n12090), .D(n12810), .Z(n5_adj_7936)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_3_lut_4_lut_adj_171.init = 16'h6996;
    LUT4 i2_2_lut_3_lut_4_lut_adj_172 (.A(block_new_127__N_1901[118]), .B(block_new_127__N_1901[108]), 
         .C(block_new_127__N_1901[102]), .D(block_new_127__N_1901[110]), 
         .Z(n7_adj_7883)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i2_2_lut_3_lut_4_lut_adj_172.init = 16'h6996;
    LUT4 i3_3_lut_4_lut_adj_173 (.A(block_new_127__N_1901[118]), .B(block_new_127__N_1901[108]), 
         .C(n33836), .D(n33831), .Z(n8_adj_8001)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i3_3_lut_4_lut_adj_173.init = 16'h6996;
    LUT4 i2_3_lut_rep_487 (.A(block_new_127__N_1901[125]), .B(block_new_127__N_1901[101]), 
         .C(block_new_127__N_1901[117]), .Z(n33791)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i2_3_lut_rep_487.init = 16'h9696;
    LUT4 i1_2_lut_rep_375_4_lut (.A(block_new_127__N_1901[125]), .B(block_new_127__N_1901[101]), 
         .C(block_new_127__N_1901[117]), .D(block_new_127__N_1901[109]), 
         .Z(n33679)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_375_4_lut.init = 16'h6996;
    LUT4 i2_2_lut_3_lut_4_lut_adj_174 (.A(block_new_127__N_1901[75]), .B(block_new_127__N_1901[79]), 
         .C(block_new_127__N_1901[68]), .D(n12748), .Z(n6_adj_7897)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i2_2_lut_3_lut_4_lut_adj_174.init = 16'h6996;
    LUT4 i1_2_lut_rep_379_3_lut_4_lut (.A(block_new_127__N_1901[91]), .B(block_new_127__N_1901[95]), 
         .C(block_new_127__N_1901[79]), .D(block_new_127__N_1901[75]), .Z(n33683)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_379_3_lut_4_lut.init = 16'h6996;
    LUT4 i2_2_lut_3_lut_4_lut_adj_175 (.A(block_new_127__N_1901[91]), .B(block_new_127__N_1901[95]), 
         .C(n33705), .D(n33797), .Z(n7_adj_7949)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i2_2_lut_3_lut_4_lut_adj_175.init = 16'h6996;
    LUT4 i3_3_lut_4_lut_adj_176 (.A(block_new_127__N_1901[84]), .B(block_new_127__N_1901[92]), 
         .C(n12748), .D(block_new_127__N_1901[76]), .Z(n8_adj_7950)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i3_3_lut_4_lut_adj_176.init = 16'h6996;
    LUT4 i2_3_lut_rep_277_4_lut (.A(block_new_127__N_1901[97]), .B(n33768), 
         .C(block_new_127__N_1901[110]), .D(block_new_127__N_1901[105]), 
         .Z(n33581)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i2_3_lut_rep_277_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_399_3_lut (.A(block_new_127__N_1901[83]), .B(block_new_127__N_1901[87]), 
         .C(block_new_127__N_1901[68]), .Z(n33703)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_399_3_lut.init = 16'h9696;
    LUT4 i1_2_lut_rep_284_3_lut_4_lut (.A(block_new_127__N_1901[83]), .B(block_new_127__N_1901[87]), 
         .C(block_new_127__N_1901[85]), .D(block_new_127__N_1901[68]), .Z(n33588)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_284_3_lut_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_398_3_lut (.A(block_new_127__N_1901[83]), .B(block_new_127__N_1901[87]), 
         .C(block_new_127__N_1901[76]), .Z(n33702)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_398_3_lut.init = 16'h9696;
    LUT4 i1_2_lut_3_lut_4_lut_adj_177 (.A(block_new_127__N_1901[83]), .B(block_new_127__N_1901[87]), 
         .C(block_new_127__N_1901[68]), .D(block_new_127__N_1901[76]), .Z(n5_adj_7926)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_3_lut_4_lut_adj_177.init = 16'h6996;
    LUT4 i1_2_lut_rep_377_3_lut (.A(block_new_127__N_1901[78]), .B(block_new_127__N_1901[94]), 
         .C(block_new_127__N_1901[77]), .Z(n33681)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_rep_377_3_lut.init = 16'h9696;
    LUT4 i1_2_lut_4_lut_adj_178 (.A(block_new_127__N_1901[72]), .B(n33804), 
         .C(block_new_127__N_1901[95]), .D(block_new_127__N_1901[80]), .Z(n5_adj_7761)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_4_lut_adj_178.init = 16'h6996;
    LUT4 block_127__I_0_i128_2_lut (.A(\block_reg[0] [31]), .B(round_key[127]), 
         .Z(block_new_127__N_1645_c[127])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i128_2_lut.init = 16'h6666;
    LUT4 i2_3_lut_rep_400_4_lut (.A(block_new_127__N_1901[78]), .B(block_new_127__N_1901[94]), 
         .C(n33809), .D(n33822), .Z(n33704)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i2_3_lut_rep_400_4_lut.init = 16'h6996;
    FD1P3AX block_w3_reg__i2 (.D(n3899[1]), .SP(block_w3_we), .CK(clk_c), 
            .Q(dec_new_block[1])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w3_reg__i2.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i3 (.D(n3899[2]), .SP(block_w3_we), .CK(clk_c), 
            .Q(dec_new_block[2])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w3_reg__i3.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i4 (.D(n3899[3]), .SP(block_w3_we), .CK(clk_c), 
            .Q(dec_new_block[3])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w3_reg__i4.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i5 (.D(n3899[4]), .SP(block_w3_we), .CK(clk_c), 
            .Q(dec_new_block[4])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w3_reg__i5.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i6 (.D(n3899[5]), .SP(block_w3_we), .CK(clk_c), 
            .Q(dec_new_block[5])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w3_reg__i6.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i7 (.D(n3899[6]), .SP(block_w3_we), .CK(clk_c), 
            .Q(dec_new_block[6])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w3_reg__i7.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i8 (.D(n3899[7]), .SP(block_w3_we), .CK(clk_c), 
            .Q(dec_new_block[7])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w3_reg__i8.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i9 (.D(n3899[8]), .SP(block_w3_we), .CK(clk_c), 
            .Q(dec_new_block[8])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w3_reg__i9.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i10 (.D(n3899[9]), .SP(block_w3_we), .CK(clk_c), 
            .Q(dec_new_block[9])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w3_reg__i10.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i11 (.D(n3899[10]), .SP(block_w3_we), .CK(clk_c), 
            .Q(dec_new_block[10])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w3_reg__i11.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i12 (.D(n3899[11]), .SP(block_w3_we), .CK(clk_c), 
            .Q(dec_new_block[11])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w3_reg__i12.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i13 (.D(n3899[12]), .SP(block_w3_we), .CK(clk_c), 
            .Q(dec_new_block[12])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w3_reg__i13.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i14 (.D(n3899[13]), .SP(block_w3_we), .CK(clk_c), 
            .Q(dec_new_block[13])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w3_reg__i14.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i15 (.D(n3899[14]), .SP(block_w3_we), .CK(clk_c), 
            .Q(dec_new_block[14])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w3_reg__i15.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i16 (.D(n3899[15]), .SP(block_w3_we), .CK(clk_c), 
            .Q(dec_new_block[15])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w3_reg__i16.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i17 (.D(n3899[16]), .SP(block_w3_we), .CK(clk_c), 
            .Q(dec_new_block[16])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w3_reg__i17.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i18 (.D(n3899[17]), .SP(block_w3_we), .CK(clk_c), 
            .Q(dec_new_block[17])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w3_reg__i18.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i19 (.D(n3899[18]), .SP(block_w3_we), .CK(clk_c), 
            .Q(dec_new_block[18])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w3_reg__i19.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i20 (.D(n3899[19]), .SP(block_w3_we), .CK(clk_c), 
            .Q(dec_new_block[19])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w3_reg__i20.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i21 (.D(n3899[20]), .SP(block_w3_we), .CK(clk_c), 
            .Q(dec_new_block[20])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w3_reg__i21.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i22 (.D(n3899[21]), .SP(block_w3_we), .CK(clk_c), 
            .Q(dec_new_block[21])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w3_reg__i22.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i23 (.D(n3899[22]), .SP(block_w3_we), .CK(clk_c), 
            .Q(dec_new_block[22])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w3_reg__i23.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i24 (.D(n3899[23]), .SP(block_w3_we), .CK(clk_c), 
            .Q(dec_new_block[23])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w3_reg__i24.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i25 (.D(n3899[24]), .SP(block_w3_we), .CK(clk_c), 
            .Q(dec_new_block[24])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w3_reg__i25.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i26 (.D(n3899[25]), .SP(block_w3_we), .CK(clk_c), 
            .Q(dec_new_block[25])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w3_reg__i26.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i27 (.D(n3899[26]), .SP(block_w3_we), .CK(clk_c), 
            .Q(dec_new_block[26])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w3_reg__i27.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i28 (.D(n3899[27]), .SP(block_w3_we), .CK(clk_c), 
            .Q(dec_new_block[27])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w3_reg__i28.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i29 (.D(n3899[28]), .SP(block_w3_we), .CK(clk_c), 
            .Q(dec_new_block[28])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w3_reg__i29.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i30 (.D(n3899[29]), .SP(block_w3_we), .CK(clk_c), 
            .Q(dec_new_block[29])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w3_reg__i30.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i31 (.D(n3899[30]), .SP(block_w3_we), .CK(clk_c), 
            .Q(dec_new_block[30])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w3_reg__i31.GSR = "ENABLED";
    FD1P3AX block_w3_reg__i32 (.D(n3899[31]), .SP(block_w3_we), .CK(clk_c), 
            .Q(dec_new_block[31])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w3_reg__i32.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_179 (.A(dec_ctrl_new_2__N_2032), .B(n6363[1]), .C(n6363[2]), 
         .D(n33856), .Z(update_type[0])) /* synthesis lut_function=(!(A+!(B (C)+!B (C+(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(197[17:30])
    defparam i1_4_lut_adj_179.init = 16'h5150;
    LUT4 block_127__I_0_i127_2_lut (.A(\block_reg[0] [30]), .B(round_key[126]), 
         .Z(block_new_127__N_1645_c[126])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i127_2_lut.init = 16'h6666;
    LUT4 i4_4_lut (.A(n33812), .B(n33748), .C(block_new_127__N_1901[53]), 
         .D(n33764), .Z(n10_adj_8002)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i4_4_lut.init = 16'h6996;
    FD1P3AX round_ctr_reg_i0_i1 (.D(round_ctr_new_c[1]), .SP(round_ctr_we), 
            .CK(clk_c), .Q(dec_round_nr_c[1])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam round_ctr_reg_i0_i1.GSR = "ENABLED";
    FD1P3AX round_ctr_reg_i0_i2 (.D(round_ctr_new_c[2]), .SP(round_ctr_we), 
            .CK(clk_c), .Q(dec_round_nr_c[2])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam round_ctr_reg_i0_i2.GSR = "ENABLED";
    FD1P3AX round_ctr_reg_i0_i3 (.D(\round_ctr_new[3] ), .SP(round_ctr_we), 
            .CK(clk_c), .Q(dec_round_nr_c[3])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam round_ctr_reg_i0_i3.GSR = "ENABLED";
    LUT4 i5_4_lut (.A(block_new_127__N_1901[127]), .B(block_new_127__N_1901[102]), 
         .C(n12084), .D(block_new_127__N_1901[124]), .Z(n12_adj_8003)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i5_4_lut.init = 16'h6996;
    LUT4 i3_3_lut_4_lut_adj_180 (.A(block_new_127__N_1901[77]), .B(n33795), 
         .C(n33680), .D(block_new_127__N_1901[93]), .Z(n8_adj_7851)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i3_3_lut_4_lut_adj_180.init = 16'h6996;
    LUT4 i3_3_lut_rep_401_4_lut (.A(block_new_127__N_1901[70]), .B(block_new_127__N_1901[86]), 
         .C(n33821), .D(n33816), .Z(n33705)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i3_3_lut_rep_401_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_273_3_lut_4_lut (.A(block_new_127__N_1901[70]), .B(block_new_127__N_1901[86]), 
         .C(n33803), .D(block_new_127__N_1901[88]), .Z(n33577)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_rep_273_3_lut_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_536_4_lut (.A(dec_new_block[126]), .B(round_key[126]), 
         .C(dec_new_block[111]), .D(round_key[111]), .Z(n33840)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_536_4_lut.init = 16'h6996;
    LUT4 xor_54_i5_2_lut_rep_534_4_lut (.A(dec_new_block[107]), .B(round_key[107]), 
         .C(dec_new_block[111]), .D(round_key[111]), .Z(n33838)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam xor_54_i5_2_lut_rep_534_4_lut.init = 16'h6996;
    LUT4 xor_29_i5_2_lut_rep_533_4_lut (.A(dec_new_block[123]), .B(round_key[123]), 
         .C(dec_new_block[127]), .D(round_key[127]), .Z(n33837)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam xor_29_i5_2_lut_rep_533_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_3_lut_adj_181 (.A(block_new_127__N_1901[67]), .B(block_new_127__N_1901[71]), 
         .C(block_new_127__N_1901[84]), .Z(n29381)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_3_lut_adj_181.init = 16'h9696;
    FD1P3AX block_w1_reg__i2 (.D(n3899[65]), .SP(block_w1_we), .CK(clk_c), 
            .Q(dec_new_block[65])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w1_reg__i2.GSR = "ENABLED";
    LUT4 mux_626_Mux_23_i2_4_lut (.A(new_sboxw[23]), .B(n33576), .C(update_type[0]), 
         .D(n4_adj_7998), .Z(n2_adj_8004)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_23_i2_4_lut.init = 16'h3aca;
    FD1P3AX block_w1_reg__i3 (.D(n3899[66]), .SP(block_w1_we), .CK(clk_c), 
            .Q(dec_new_block[66])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w1_reg__i3.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i4 (.D(n3899[67]), .SP(block_w1_we), .CK(clk_c), 
            .Q(dec_new_block[67])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w1_reg__i4.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i5 (.D(n3899[68]), .SP(block_w1_we), .CK(clk_c), 
            .Q(dec_new_block[68])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w1_reg__i5.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i6 (.D(n3899[69]), .SP(block_w1_we), .CK(clk_c), 
            .Q(dec_new_block[69])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w1_reg__i6.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i7 (.D(n3899[70]), .SP(block_w1_we), .CK(clk_c), 
            .Q(dec_new_block[70])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w1_reg__i7.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i8 (.D(n3899[71]), .SP(block_w1_we), .CK(clk_c), 
            .Q(dec_new_block[71])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w1_reg__i8.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i9 (.D(n3899[72]), .SP(block_w1_we), .CK(clk_c), 
            .Q(dec_new_block[72])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w1_reg__i9.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i10 (.D(n3899[73]), .SP(block_w1_we), .CK(clk_c), 
            .Q(dec_new_block[73])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w1_reg__i10.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i11 (.D(n3899[74]), .SP(block_w1_we), .CK(clk_c), 
            .Q(dec_new_block[74])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w1_reg__i11.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i12 (.D(n3899[75]), .SP(block_w1_we), .CK(clk_c), 
            .Q(dec_new_block[75])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w1_reg__i12.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i13 (.D(n3899[76]), .SP(block_w1_we), .CK(clk_c), 
            .Q(dec_new_block[76])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w1_reg__i13.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i14 (.D(n3899[77]), .SP(block_w1_we), .CK(clk_c), 
            .Q(dec_new_block[77])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w1_reg__i14.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i15 (.D(n3899[78]), .SP(block_w1_we), .CK(clk_c), 
            .Q(dec_new_block[78])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w1_reg__i15.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i16 (.D(n3899[79]), .SP(block_w1_we), .CK(clk_c), 
            .Q(dec_new_block[79])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w1_reg__i16.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i17 (.D(n3899[80]), .SP(block_w1_we), .CK(clk_c), 
            .Q(dec_new_block[80])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w1_reg__i17.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i18 (.D(n3899[81]), .SP(block_w1_we), .CK(clk_c), 
            .Q(dec_new_block[81])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w1_reg__i18.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i19 (.D(n3899[82]), .SP(block_w1_we), .CK(clk_c), 
            .Q(dec_new_block[82])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w1_reg__i19.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i20 (.D(n3899[83]), .SP(block_w1_we), .CK(clk_c), 
            .Q(dec_new_block[83])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w1_reg__i20.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i21 (.D(n3899[84]), .SP(block_w1_we), .CK(clk_c), 
            .Q(dec_new_block[84])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w1_reg__i21.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i22 (.D(n3899[85]), .SP(block_w1_we), .CK(clk_c), 
            .Q(dec_new_block[85])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w1_reg__i22.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i23 (.D(n3899[86]), .SP(block_w1_we), .CK(clk_c), 
            .Q(dec_new_block[86])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w1_reg__i23.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i24 (.D(n3899[87]), .SP(block_w1_we), .CK(clk_c), 
            .Q(dec_new_block[87])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w1_reg__i24.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i25 (.D(n3899[88]), .SP(block_w1_we), .CK(clk_c), 
            .Q(dec_new_block[88])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w1_reg__i25.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i26 (.D(n3899[89]), .SP(block_w1_we), .CK(clk_c), 
            .Q(dec_new_block[89])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w1_reg__i26.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i27 (.D(n3899[90]), .SP(block_w1_we), .CK(clk_c), 
            .Q(dec_new_block[90])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w1_reg__i27.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i28 (.D(n3899[91]), .SP(block_w1_we), .CK(clk_c), 
            .Q(dec_new_block[91])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w1_reg__i28.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i29 (.D(n3899[92]), .SP(block_w1_we), .CK(clk_c), 
            .Q(dec_new_block[92])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w1_reg__i29.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i30 (.D(n3899[93]), .SP(block_w1_we), .CK(clk_c), 
            .Q(dec_new_block[93])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w1_reg__i30.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i31 (.D(n3899[94]), .SP(block_w1_we), .CK(clk_c), 
            .Q(dec_new_block[94])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w1_reg__i31.GSR = "ENABLED";
    FD1P3AX block_w1_reg__i32 (.D(n3899[95]), .SP(block_w1_we), .CK(clk_c), 
            .Q(dec_new_block[95])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w1_reg__i32.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i2 (.D(n3899[97]), .SP(block_w0_we), .CK(clk_c), 
            .Q(dec_new_block[97])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w0_reg__i2.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i3 (.D(n3899[98]), .SP(block_w0_we), .CK(clk_c), 
            .Q(dec_new_block[98])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w0_reg__i3.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i4 (.D(n3899[99]), .SP(block_w0_we), .CK(clk_c), 
            .Q(dec_new_block[99])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w0_reg__i4.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i5 (.D(n3899[100]), .SP(block_w0_we), .CK(clk_c), 
            .Q(dec_new_block[100])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w0_reg__i5.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i6 (.D(n3899[101]), .SP(block_w0_we), .CK(clk_c), 
            .Q(dec_new_block[101])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w0_reg__i6.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i7 (.D(n3899[102]), .SP(block_w0_we), .CK(clk_c), 
            .Q(dec_new_block[102])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w0_reg__i7.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i8 (.D(n3899[103]), .SP(block_w0_we), .CK(clk_c), 
            .Q(dec_new_block[103])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w0_reg__i8.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i9 (.D(n3899[104]), .SP(block_w0_we), .CK(clk_c), 
            .Q(dec_new_block[104])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w0_reg__i9.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i10 (.D(n3899[105]), .SP(block_w0_we), .CK(clk_c), 
            .Q(dec_new_block[105])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w0_reg__i10.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i11 (.D(n3899[106]), .SP(block_w0_we), .CK(clk_c), 
            .Q(dec_new_block[106])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w0_reg__i11.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i12 (.D(n3899[107]), .SP(block_w0_we), .CK(clk_c), 
            .Q(dec_new_block[107])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w0_reg__i12.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i13 (.D(n3899[108]), .SP(block_w0_we), .CK(clk_c), 
            .Q(dec_new_block[108])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w0_reg__i13.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i14 (.D(n3899[109]), .SP(block_w0_we), .CK(clk_c), 
            .Q(dec_new_block[109])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w0_reg__i14.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i15 (.D(n3899[110]), .SP(block_w0_we), .CK(clk_c), 
            .Q(dec_new_block[110])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w0_reg__i15.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i16 (.D(n3899[111]), .SP(block_w0_we), .CK(clk_c), 
            .Q(dec_new_block[111])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w0_reg__i16.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i17 (.D(n3899[112]), .SP(block_w0_we), .CK(clk_c), 
            .Q(dec_new_block[112])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w0_reg__i17.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i18 (.D(n3899[113]), .SP(block_w0_we), .CK(clk_c), 
            .Q(dec_new_block[113])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w0_reg__i18.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i19 (.D(n3899[114]), .SP(block_w0_we), .CK(clk_c), 
            .Q(dec_new_block[114])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w0_reg__i19.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i20 (.D(n3899[115]), .SP(block_w0_we), .CK(clk_c), 
            .Q(dec_new_block[115])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w0_reg__i20.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i21 (.D(n3899[116]), .SP(block_w0_we), .CK(clk_c), 
            .Q(dec_new_block[116])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w0_reg__i21.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i22 (.D(n3899[117]), .SP(block_w0_we), .CK(clk_c), 
            .Q(dec_new_block[117])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w0_reg__i22.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i23 (.D(n3899[118]), .SP(block_w0_we), .CK(clk_c), 
            .Q(dec_new_block[118])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w0_reg__i23.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i24 (.D(n3899[119]), .SP(block_w0_we), .CK(clk_c), 
            .Q(dec_new_block[119])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w0_reg__i24.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i25 (.D(n3899[120]), .SP(block_w0_we), .CK(clk_c), 
            .Q(dec_new_block[120])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w0_reg__i25.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i26 (.D(n3899[121]), .SP(block_w0_we), .CK(clk_c), 
            .Q(dec_new_block[121])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w0_reg__i26.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i27 (.D(n3899[122]), .SP(block_w0_we), .CK(clk_c), 
            .Q(dec_new_block[122])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w0_reg__i27.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i28 (.D(n3899[123]), .SP(block_w0_we), .CK(clk_c), 
            .Q(dec_new_block[123])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w0_reg__i28.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i29 (.D(n3899[124]), .SP(block_w0_we), .CK(clk_c), 
            .Q(dec_new_block[124])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w0_reg__i29.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i30 (.D(n3899[125]), .SP(block_w0_we), .CK(clk_c), 
            .Q(dec_new_block[125])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w0_reg__i30.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i31 (.D(n3899[126]), .SP(block_w0_we), .CK(clk_c), 
            .Q(dec_new_block[126])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w0_reg__i31.GSR = "ENABLED";
    FD1P3AX block_w0_reg__i32 (.D(n3899[127]), .SP(block_w0_we), .CK(clk_c), 
            .Q(dec_new_block[127])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w0_reg__i32.GSR = "ENABLED";
    LUT4 i2_2_lut_4_lut_adj_182 (.A(dec_new_block[95]), .B(round_key[95]), 
         .C(dec_new_block[70]), .D(round_key[70]), .Z(n7_adj_7700)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i2_2_lut_4_lut_adj_182.init = 16'h6996;
    LUT4 i2_2_lut_4_lut_adj_183 (.A(dec_new_block[7]), .B(round_key[7]), 
         .C(dec_new_block[16]), .D(round_key[16]), .Z(n7_adj_7709)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i2_2_lut_4_lut_adj_183.init = 16'h6996;
    LUT4 i1_2_lut_rep_532_4_lut (.A(dec_new_block[117]), .B(round_key[117]), 
         .C(dec_new_block[124]), .D(round_key[124]), .Z(n33836)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_rep_532_4_lut.init = 16'h6996;
    LUT4 i1_4_lut_adj_184 (.A(encdec_reg), .B(n14890), .C(dec_ready), 
         .D(n33942), .Z(n6431)) /* synthesis lut_function=(A (B+(C))+!A (B+!((D)+!C))) */ ;
    defparam i1_4_lut_adj_184.init = 16'hecfc;
    LUT4 xor_43_i4_2_lut_rep_531_4_lut (.A(dec_new_block[114]), .B(round_key[114]), 
         .C(dec_new_block[119]), .D(round_key[119]), .Z(n33835)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam xor_43_i4_2_lut_rep_531_4_lut.init = 16'h6996;
    FD1P3AX block_w2_reg__i2 (.D(n3899[33]), .SP(block_w2_we), .CK(clk_c), 
            .Q(dec_new_block[33])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w2_reg__i2.GSR = "ENABLED";
    LUT4 new_block_127__I_0_i120_2_lut (.A(dec_new_block[119]), .B(round_key[119]), 
         .Z(block_new_127__N_1901[119])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i120_2_lut.init = 16'h6666;
    LUT4 i1_2_lut_rep_388_3_lut (.A(block_new_127__N_1901[67]), .B(block_new_127__N_1901[71]), 
         .C(block_new_127__N_1901[92]), .Z(n33692)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_388_3_lut.init = 16'h9696;
    LUT4 i1_2_lut_rep_394_3_lut (.A(block_new_127__N_1901[43]), .B(block_new_127__N_1901[47]), 
         .C(block_new_127__N_1901[37]), .Z(n33698)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_394_3_lut.init = 16'h9696;
    LUT4 i2_2_lut_3_lut_adj_185 (.A(block_new_127__N_1901[43]), .B(block_new_127__N_1901[47]), 
         .C(block_new_127__N_1901[61]), .Z(n7_adj_7862)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i2_2_lut_3_lut_adj_185.init = 16'h9696;
    LUT4 i3_3_lut_4_lut_adj_186 (.A(block_new_127__N_1901[77]), .B(n33795), 
         .C(block_new_127__N_1901[70]), .D(n29381), .Z(n8_adj_7725)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i3_3_lut_4_lut_adj_186.init = 16'h6996;
    LUT4 i1_2_lut_rep_403_3_lut_4_lut (.A(block_new_127__N_1901[35]), .B(block_new_127__N_1901[39]), 
         .C(block_new_127__N_1901[47]), .D(block_new_127__N_1901[43]), .Z(n33707)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_403_3_lut_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_3_lut_adj_187 (.A(block_new_127__N_1901[60]), .B(block_new_127__N_1901[52]), 
         .C(block_new_127__N_1901[36]), .Z(n5_adj_7955)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_3_lut_adj_187.init = 16'h9696;
    LUT4 i1_2_lut_3_lut_adj_188 (.A(block_new_127__N_1901[60]), .B(block_new_127__N_1901[52]), 
         .C(n12921), .Z(n5_adj_7836)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_3_lut_adj_188.init = 16'h9696;
    LUT4 i1_2_lut_rep_366_3_lut (.A(block_new_127__N_1901[62]), .B(block_new_127__N_1901[46]), 
         .C(block_new_127__N_1901[53]), .Z(n33670)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_rep_366_3_lut.init = 16'h9696;
    LUT4 i2_3_lut_rep_402_4_lut (.A(block_new_127__N_1901[62]), .B(block_new_127__N_1901[46]), 
         .C(n33814), .D(n33805), .Z(n33706)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i2_3_lut_rep_402_4_lut.init = 16'h6996;
    LUT4 i2_2_lut_3_lut_adj_189 (.A(block_new_127__N_1901[53]), .B(block_new_127__N_1901[61]), 
         .C(n29408), .Z(n7_adj_8005)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i2_2_lut_3_lut_adj_189.init = 16'h9696;
    LUT4 i2_2_lut_4_lut_adj_190 (.A(n33711), .B(block_new_127__N_1901[33]), 
         .C(n12071), .D(n33760), .Z(n6_adj_7703)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i2_2_lut_4_lut_adj_190.init = 16'h6996;
    FD1P3AX block_w2_reg__i3 (.D(n3899[34]), .SP(block_w2_we), .CK(clk_c), 
            .Q(dec_new_block[34])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w2_reg__i3.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i4 (.D(n3899[35]), .SP(block_w2_we), .CK(clk_c), 
            .Q(dec_new_block[35])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w2_reg__i4.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i5 (.D(n3899[36]), .SP(block_w2_we), .CK(clk_c), 
            .Q(dec_new_block[36])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w2_reg__i5.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i6 (.D(n3899[37]), .SP(block_w2_we), .CK(clk_c), 
            .Q(dec_new_block[37])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w2_reg__i6.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i7 (.D(n3899[38]), .SP(block_w2_we), .CK(clk_c), 
            .Q(dec_new_block[38])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w2_reg__i7.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i8 (.D(n3899[39]), .SP(block_w2_we), .CK(clk_c), 
            .Q(dec_new_block[39])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w2_reg__i8.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i9 (.D(n3899[40]), .SP(block_w2_we), .CK(clk_c), 
            .Q(dec_new_block[40])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w2_reg__i9.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i10 (.D(n3899[41]), .SP(block_w2_we), .CK(clk_c), 
            .Q(dec_new_block[41])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w2_reg__i10.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i11 (.D(n3899[42]), .SP(block_w2_we), .CK(clk_c), 
            .Q(dec_new_block[42])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w2_reg__i11.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i12 (.D(n3899[43]), .SP(block_w2_we), .CK(clk_c), 
            .Q(dec_new_block[43])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w2_reg__i12.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i13 (.D(n3899[44]), .SP(block_w2_we), .CK(clk_c), 
            .Q(dec_new_block[44])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w2_reg__i13.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i14 (.D(n3899[45]), .SP(block_w2_we), .CK(clk_c), 
            .Q(dec_new_block[45])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w2_reg__i14.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i15 (.D(n3899[46]), .SP(block_w2_we), .CK(clk_c), 
            .Q(dec_new_block[46])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w2_reg__i15.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i16 (.D(n3899[47]), .SP(block_w2_we), .CK(clk_c), 
            .Q(dec_new_block[47])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w2_reg__i16.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i17 (.D(n3899[48]), .SP(block_w2_we), .CK(clk_c), 
            .Q(dec_new_block[48])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w2_reg__i17.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i18 (.D(n3899[49]), .SP(block_w2_we), .CK(clk_c), 
            .Q(dec_new_block[49])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w2_reg__i18.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i19 (.D(n3899[50]), .SP(block_w2_we), .CK(clk_c), 
            .Q(dec_new_block[50])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w2_reg__i19.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i20 (.D(n3899[51]), .SP(block_w2_we), .CK(clk_c), 
            .Q(dec_new_block[51])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w2_reg__i20.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i21 (.D(n3899[52]), .SP(block_w2_we), .CK(clk_c), 
            .Q(dec_new_block[52])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w2_reg__i21.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i22 (.D(n3899[53]), .SP(block_w2_we), .CK(clk_c), 
            .Q(dec_new_block[53])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w2_reg__i22.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i23 (.D(n3899[54]), .SP(block_w2_we), .CK(clk_c), 
            .Q(dec_new_block[54])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w2_reg__i23.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i24 (.D(n3899[55]), .SP(block_w2_we), .CK(clk_c), 
            .Q(dec_new_block[55])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w2_reg__i24.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i25 (.D(n3899[56]), .SP(block_w2_we), .CK(clk_c), 
            .Q(dec_new_block[56])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w2_reg__i25.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i26 (.D(n3899[57]), .SP(block_w2_we), .CK(clk_c), 
            .Q(dec_new_block[57])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w2_reg__i26.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i27 (.D(n3899[58]), .SP(block_w2_we), .CK(clk_c), 
            .Q(dec_new_block[58])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w2_reg__i27.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i28 (.D(n3899[59]), .SP(block_w2_we), .CK(clk_c), 
            .Q(dec_new_block[59])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w2_reg__i28.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i29 (.D(n3899[60]), .SP(block_w2_we), .CK(clk_c), 
            .Q(dec_new_block[60])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w2_reg__i29.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i30 (.D(n3899[61]), .SP(block_w2_we), .CK(clk_c), 
            .Q(dec_new_block[61])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w2_reg__i30.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i31 (.D(n3899[62]), .SP(block_w2_we), .CK(clk_c), 
            .Q(dec_new_block[62])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w2_reg__i31.GSR = "ENABLED";
    FD1P3AX block_w2_reg__i32 (.D(n3899[63]), .SP(block_w2_we), .CK(clk_c), 
            .Q(dec_new_block[63])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=22, LSE_RCOL=32, LSE_LLINE=135, LSE_RLINE=148 */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(268[9] 292[12])
    defparam block_w2_reg__i32.GSR = "ENABLED";
    LUT4 mux_626_Mux_48_i2_4_lut (.A(new_sboxw[16]), .B(n33577), .C(update_type[0]), 
         .D(n4_adj_7680), .Z(n2_adj_8006)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_48_i2_4_lut.init = 16'h3aca;
    LUT4 n2753_bdd_4_lut (.A(n2752[31]), .B(n9426), .C(n30146), .D(n25333), 
         .Z(tmp_sboxw[31])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n2753_bdd_4_lut.init = 16'h00ca;
    LUT4 xor_67_i4_2_lut_rep_530_4_lut (.A(dec_new_block[98]), .B(round_key[98]), 
         .C(dec_new_block[103]), .D(round_key[103]), .Z(n33834)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam xor_67_i4_2_lut_rep_530_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_4_lut_adj_191 (.A(dec_new_block[119]), .B(round_key[119]), 
         .C(dec_new_block[104]), .D(round_key[104]), .Z(n5_adj_7780)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_4_lut_adj_191.init = 16'h6996;
    LUT4 xor_54_i4_2_lut_rep_529_4_lut (.A(dec_new_block[106]), .B(round_key[106]), 
         .C(dec_new_block[111]), .D(round_key[111]), .Z(n33833)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam xor_54_i4_2_lut_rep_529_4_lut.init = 16'h6996;
    LUT4 i2_3_lut_rep_271_4_lut (.A(block_new_127__N_1901[37]), .B(n33812), 
         .C(n12071), .D(block_new_127__N_1901[33]), .Z(n33575)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i2_3_lut_rep_271_4_lut.init = 16'h6996;
    LUT4 mux_626_Mux_55_i2_4_lut (.A(new_sboxw[23]), .B(n33578), .C(update_type[0]), 
         .D(n4_adj_7813), .Z(n2_adj_8007)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_55_i2_4_lut.init = 16'h3aca;
    LUT4 i1_2_lut_4_lut_adj_192 (.A(dec_new_block[97]), .B(round_key[97]), 
         .C(dec_new_block[122]), .D(round_key[122]), .Z(n5_adj_7785)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_4_lut_adj_192.init = 16'h6996;
    LUT4 xor_29_i4_2_lut_rep_528_4_lut (.A(dec_new_block[122]), .B(round_key[122]), 
         .C(dec_new_block[127]), .D(round_key[127]), .Z(n33832)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam xor_29_i4_2_lut_rep_528_4_lut.init = 16'h6996;
    LUT4 i2_2_lut_3_lut_adj_193 (.A(dec_new_block[81]), .B(round_key[81]), 
         .C(n29146), .Z(n6_adj_7854)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i2_2_lut_3_lut_adj_193.init = 16'h9696;
    LUT4 i1_2_lut_rep_527_4_lut (.A(dec_new_block[101]), .B(round_key[101]), 
         .C(dec_new_block[103]), .D(round_key[103]), .Z(n33831)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_527_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_3_lut_4_lut_adj_194 (.A(block_new_127__N_1901[37]), .B(n33812), 
         .C(n33787), .D(block_new_127__N_1901[52]), .Z(n5_adj_7803)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_3_lut_4_lut_adj_194.init = 16'h6996;
    LUT4 i2_2_lut_3_lut_adj_195 (.A(dec_new_block[4]), .B(round_key[4]), 
         .C(n29143), .Z(n7_adj_7874)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i2_2_lut_3_lut_adj_195.init = 16'h9696;
    LUT4 mux_626_Mux_58_i2_4_lut (.A(new_sboxw[26]), .B(n5_adj_7752), .C(update_type[0]), 
         .D(n6_adj_8008), .Z(n2_adj_8009)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_58_i2_4_lut.init = 16'h3aca;
    LUT4 i2_2_lut_4_lut_adj_196 (.A(dec_new_block[98]), .B(round_key[98]), 
         .C(dec_new_block[110]), .D(round_key[110]), .Z(n7_adj_7877)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i2_2_lut_4_lut_adj_196.init = 16'h6996;
    LUT4 i1_2_lut_4_lut_adj_197 (.A(dec_new_block[125]), .B(round_key[125]), 
         .C(dec_new_block[118]), .D(round_key[118]), .Z(n5_adj_7885)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_4_lut_adj_197.init = 16'h6996;
    LUT4 i1_2_lut_rep_526_4_lut (.A(dec_new_block[109]), .B(round_key[109]), 
         .C(dec_new_block[111]), .D(round_key[111]), .Z(n33830)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_526_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_3_lut_adj_198 (.A(dec_new_block[32]), .B(round_key[32]), 
         .C(n28926), .Z(n4_adj_7899)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_3_lut_adj_198.init = 16'h9696;
    LUT4 i1_2_lut_3_lut_adj_199 (.A(dec_new_block[10]), .B(round_key[10]), 
         .C(n28882), .Z(n4_adj_7905)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_3_lut_adj_199.init = 16'h9696;
    LUT4 block_127__I_0_i23_2_lut (.A(\block_reg[3] [22]), .B(round_key[22]), 
         .Z(block_new_127__N_1645_c[22])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i23_2_lut.init = 16'h6666;
    LUT4 i1_2_lut_rep_404_3_lut (.A(block_new_127__N_1901[93]), .B(block_new_127__N_1901[77]), 
         .C(block_new_127__N_1901[71]), .Z(n33708)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_rep_404_3_lut.init = 16'h9696;
    LUT4 i2_2_lut_3_lut_4_lut_adj_200 (.A(n33792), .B(n33793), .C(n33705), 
         .D(block_new_127__N_1901[93]), .Z(n6_adj_7697)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i2_2_lut_3_lut_4_lut_adj_200.init = 16'h6996;
    LUT4 i1_2_lut_3_lut_4_lut_adj_201 (.A(n33792), .B(n33793), .C(block_new_127__N_1901[78]), 
         .D(block_new_127__N_1901[93]), .Z(n5_adj_7856)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_3_lut_4_lut_adj_201.init = 16'h6996;
    LUT4 i2_3_lut_rep_217_4_lut (.A(block_new_127__N_1901[69]), .B(block_new_127__N_1901[85]), 
         .C(n33590), .D(block_new_127__N_1901[78]), .Z(n33521)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i2_3_lut_rep_217_4_lut.init = 16'h6996;
    LUT4 i2_3_lut_rep_376_4_lut (.A(block_new_127__N_1901[69]), .B(block_new_127__N_1901[85]), 
         .C(block_new_127__N_1901[95]), .D(block_new_127__N_1901[72]), .Z(n33680)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i2_3_lut_rep_376_4_lut.init = 16'h6996;
    LUT4 i2_2_lut_3_lut_4_lut_adj_202 (.A(n33792), .B(n33793), .C(n33703), 
         .D(block_new_127__N_1901[85]), .Z(n7_adj_7724)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i2_2_lut_3_lut_4_lut_adj_202.init = 16'h6996;
    LUT4 i3_3_lut_4_lut_adj_203 (.A(block_new_127__N_1901[89]), .B(block_new_127__N_1901[65]), 
         .C(block_new_127__N_1901[73]), .D(block_new_127__N_1901[80]), .Z(n8_adj_7963)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i3_3_lut_4_lut_adj_203.init = 16'h6996;
    LUT4 i3_2_lut_3_lut_4_lut_adj_204 (.A(block_new_127__N_1901[89]), .B(block_new_127__N_1901[65]), 
         .C(block_new_127__N_1901[86]), .D(block_new_127__N_1901[70]), .Z(n9_adj_7791)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i3_2_lut_3_lut_4_lut_adj_204.init = 16'h6996;
    LUT4 i1_2_lut_3_lut_adj_205 (.A(block_new_127__N_1901[89]), .B(block_new_127__N_1901[65]), 
         .C(block_new_127__N_1901[82]), .Z(n4_adj_7766)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_3_lut_adj_205.init = 16'h9696;
    LUT4 new_block_127__I_0_i119_2_lut (.A(dec_new_block[118]), .B(round_key[118]), 
         .Z(block_new_127__N_1901[118])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i119_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i22_2_lut (.A(\block_reg[3] [21]), .B(round_key[21]), 
         .Z(\block_new_127__N_1645[21] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i22_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i118_2_lut (.A(dec_new_block[117]), .B(round_key[117]), 
         .Z(block_new_127__N_1901[117])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i118_2_lut.init = 16'h6666;
    LUT4 mux_626_Mux_65_i2_4_lut (.A(new_sboxw[1]), .B(n9_adj_8010), .C(update_type[0]), 
         .D(n10_adj_8002), .Z(n2_adj_8011)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_65_i2_4_lut.init = 16'h3aca;
    LUT4 xor_629_i4_2_lut_rep_525_4_lut (.A(dec_new_block[25]), .B(round_key[25]), 
         .C(dec_new_block[30]), .D(round_key[30]), .Z(n33829)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam xor_629_i4_2_lut_rep_525_4_lut.init = 16'h6996;
    LUT4 block_127__I_0_i21_2_lut (.A(\block_reg[3] [20]), .B(round_key[20]), 
         .Z(\block_new_127__N_1645[20] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i21_2_lut.init = 16'h6666;
    LUT4 xor_489_i5_2_lut_4_lut (.A(dec_new_block[59]), .B(round_key[59]), 
         .C(dec_new_block[63]), .D(round_key[63]), .Z(n4770[4])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam xor_489_i5_2_lut_4_lut.init = 16'h6996;
    LUT4 new_block_127__I_0_i117_2_lut (.A(dec_new_block[116]), .B(round_key[116]), 
         .Z(block_new_127__N_1901[116])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i117_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i20_2_lut (.A(\block_reg[3] [19]), .B(round_key[19]), 
         .Z(\block_new_127__N_1645[19] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i20_2_lut.init = 16'h6666;
    LUT4 i1_2_lut_4_lut_adj_206 (.A(dec_new_block[20]), .B(round_key[20]), 
         .C(dec_new_block[28]), .D(round_key[28]), .Z(n12090)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_4_lut_adj_206.init = 16'h6996;
    LUT4 new_block_127__I_0_i116_2_lut (.A(dec_new_block[115]), .B(round_key[115]), 
         .Z(block_new_127__N_1901[115])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i116_2_lut.init = 16'h6666;
    LUT4 i2_2_lut_3_lut_adj_207 (.A(dec_new_block[4]), .B(round_key[4]), 
         .C(n29288), .Z(n6_adj_7937)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i2_2_lut_3_lut_adj_207.init = 16'h9696;
    LUT4 block_127__I_0_i19_2_lut (.A(\block_reg[3] [18]), .B(round_key[18]), 
         .Z(block_new_127__N_1645_c[18])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i19_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i115_2_lut (.A(dec_new_block[114]), .B(round_key[114]), 
         .Z(block_new_127__N_1901[114])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i115_2_lut.init = 16'h6666;
    LUT4 i1_4_lut_adj_208 (.A(n33913), .B(n6347[0]), .C(enc_ready), .D(n33848), 
         .Z(n6428)) /* synthesis lut_function=(A (B (D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_208.init = 16'hdc50;
    LUT4 i1_2_lut_rep_524_4_lut (.A(dec_new_block[23]), .B(round_key[23]), 
         .C(dec_new_block[16]), .D(round_key[16]), .Z(n33828)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_524_4_lut.init = 16'h6996;
    LUT4 mux_626_Mux_72_i2_4_lut (.A(new_sboxw[8]), .B(n5_adj_7981), .C(update_type[0]), 
         .D(n6_adj_8012), .Z(n2_adj_8013)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_72_i2_4_lut.init = 16'h3aca;
    LUT4 i1_2_lut_rep_523_4_lut (.A(dec_new_block[21]), .B(round_key[21]), 
         .C(dec_new_block[13]), .D(round_key[13]), .Z(n33827)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_rep_523_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_522_4_lut (.A(dec_new_block[15]), .B(round_key[15]), 
         .C(dec_new_block[8]), .D(round_key[8]), .Z(n33826)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_522_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_521_4_lut (.A(dec_new_block[31]), .B(round_key[31]), 
         .C(dec_new_block[24]), .D(round_key[24]), .Z(n33825)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_521_4_lut.init = 16'h6996;
    LUT4 block_127__I_0_i18_2_lut (.A(\block_reg[3] [17]), .B(round_key[17]), 
         .Z(\block_new_127__N_1645[17] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i18_2_lut.init = 16'h6666;
    LUT4 xor_649_i4_2_lut_rep_520_4_lut (.A(dec_new_block[10]), .B(round_key[10]), 
         .C(dec_new_block[15]), .D(round_key[15]), .Z(n33824)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam xor_649_i4_2_lut_rep_520_4_lut.init = 16'h6996;
    LUT4 i2_2_lut_3_lut_adj_209 (.A(dec_new_block[108]), .B(round_key[108]), 
         .C(n29160), .Z(n7_adj_7968)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i2_2_lut_3_lut_adj_209.init = 16'h9696;
    LUT4 new_block_127__I_0_i114_2_lut (.A(dec_new_block[113]), .B(round_key[113]), 
         .Z(block_new_127__N_1901[113])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i114_2_lut.init = 16'h6666;
    LUT4 mux_626_Mux_87_i2_4_lut (.A(new_sboxw[23]), .B(n7_adj_7958), .C(update_type[0]), 
         .D(n8_adj_8001), .Z(n2_adj_8014)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_87_i2_4_lut.init = 16'h3aca;
    LUT4 i1_2_lut_rep_272_4_lut (.A(n33763), .B(block_new_127__N_1901[53]), 
         .C(block_new_127__N_1901[37]), .D(n33800), .Z(n33576)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_rep_272_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_4_lut_adj_210 (.A(n29339), .B(n33833), .C(n33832), .D(n33791), 
         .Z(n5_adj_7924)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_4_lut_adj_210.init = 16'h6996;
    LUT4 i1_4_lut_adj_211 (.A(dec_ctrl_new_2__N_2032), .B(n33842), .C(n20705), 
         .D(n33844), .Z(block_w1_we)) /* synthesis lut_function=(!(A+!(B (C+(D))+!B !((D)+!C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i1_4_lut_adj_211.init = 16'h4450;
    LUT4 mux_626_Mux_114_i2_4_lut (.A(new_sboxw[18]), .B(n7_adj_7730), .C(update_type[0]), 
         .D(n8_adj_7758), .Z(n2_adj_8015)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_114_i2_4_lut.init = 16'h3aca;
    LUT4 xor_660_i4_2_lut_rep_519_4_lut (.A(dec_new_block[2]), .B(round_key[2]), 
         .C(dec_new_block[7]), .D(round_key[7]), .Z(n33823)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam xor_660_i4_2_lut_rep_519_4_lut.init = 16'h6996;
    LUT4 xor_374_i4_2_lut_rep_518_4_lut (.A(dec_new_block[74]), .B(round_key[74]), 
         .C(dec_new_block[79]), .D(round_key[79]), .Z(n33822)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam xor_374_i4_2_lut_rep_518_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_4_lut_adj_212 (.A(dec_new_block[53]), .B(round_key[53]), 
         .C(dec_new_block[48]), .D(round_key[48]), .Z(n12071)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_4_lut_adj_212.init = 16'h6996;
    LUT4 block_127__I_0_i17_2_lut (.A(\block_reg[3] [16]), .B(round_key[16]), 
         .Z(block_new_127__N_1645_c[16])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i17_2_lut.init = 16'h6666;
    LUT4 xor_361_i4_2_lut_rep_517_4_lut (.A(dec_new_block[82]), .B(round_key[82]), 
         .C(dec_new_block[87]), .D(round_key[87]), .Z(n33821)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam xor_361_i4_2_lut_rep_517_4_lut.init = 16'h6996;
    LUT4 xor_524_i4_2_lut_4_lut (.A(dec_new_block[34]), .B(round_key[34]), 
         .C(dec_new_block[39]), .D(round_key[39]), .Z(n5085[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam xor_524_i4_2_lut_4_lut.init = 16'h6996;
    LUT4 xor_662_i4_2_lut_4_lut (.A(dec_new_block[1]), .B(round_key[1]), 
         .C(dec_new_block[6]), .D(round_key[6]), .Z(n6327[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam xor_662_i4_2_lut_4_lut.init = 16'h6996;
    LUT4 i2_2_lut_3_lut_4_lut_adj_213 (.A(n33757), .B(n33750), .C(n33779), 
         .D(n33780), .Z(n6_adj_8012)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i2_2_lut_3_lut_4_lut_adj_213.init = 16'h6996;
    LUT4 i1_2_lut_rep_516_4_lut (.A(dec_new_block[79]), .B(round_key[79]), 
         .C(dec_new_block[72]), .D(round_key[72]), .Z(n33820)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_516_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_4_lut_adj_214 (.A(dec_new_block[71]), .B(round_key[71]), 
         .C(dec_new_block[64]), .D(round_key[64]), .Z(n12074)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_4_lut_adj_214.init = 16'h6996;
    LUT4 i1_2_lut_rep_515_4_lut (.A(dec_new_block[87]), .B(round_key[87]), 
         .C(dec_new_block[80]), .D(round_key[80]), .Z(n33819)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_515_4_lut.init = 16'h6996;
    LUT4 xor_627_i4_2_lut_rep_514_4_lut (.A(dec_new_block[26]), .B(round_key[26]), 
         .C(dec_new_block[31]), .D(round_key[31]), .Z(n33818)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam xor_627_i4_2_lut_rep_514_4_lut.init = 16'h6996;
    LUT4 mux_626_Mux_119_i2_4_lut (.A(new_sboxw[23]), .B(n33574), .C(update_type[0]), 
         .D(n4_adj_7699), .Z(n2_adj_8016)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_119_i2_4_lut.init = 16'h3aca;
    LUT4 n2754_bdd_4_lut (.A(n2752[30]), .B(n9424), .C(n30146), .D(n25333), 
         .Z(tmp_sboxw[30])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n2754_bdd_4_lut.init = 16'h00ca;
    LUT4 i2_3_lut_rep_390_4_lut (.A(n29480), .B(dec_new_block[59]), .C(round_key[59]), 
         .D(block_new_127__N_1901[43]), .Z(n33694)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i2_3_lut_rep_390_4_lut.init = 16'h6996;
    LUT4 xor_634_i4_2_lut_rep_513_4_lut (.A(dec_new_block[18]), .B(round_key[18]), 
         .C(dec_new_block[23]), .D(round_key[23]), .Z(n33817)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam xor_634_i4_2_lut_rep_513_4_lut.init = 16'h6996;
    LUT4 xor_382_i4_2_lut_rep_512_4_lut (.A(dec_new_block[66]), .B(round_key[66]), 
         .C(dec_new_block[71]), .D(round_key[71]), .Z(n33816)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam xor_382_i4_2_lut_rep_512_4_lut.init = 16'h6996;
    LUT4 xor_651_i4_2_lut_4_lut (.A(dec_new_block[9]), .B(round_key[9]), 
         .C(dec_new_block[14]), .D(round_key[14]), .Z(n6228[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam xor_651_i4_2_lut_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_4_lut_adj_215 (.A(dec_new_block[112]), .B(round_key[112]), 
         .C(dec_new_block[120]), .D(round_key[120]), .Z(n29429)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_4_lut_adj_215.init = 16'h6996;
    LUT4 i4_3_lut_4_lut_adj_216 (.A(block_new_127__N_1901[101]), .B(n33839), 
         .C(block_new_127__N_1901[108]), .D(n33840), .Z(n11_adj_8017)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i4_3_lut_4_lut_adj_216.init = 16'h6996;
    LUT4 xor_56_i4_2_lut_4_lut (.A(dec_new_block[105]), .B(round_key[105]), 
         .C(dec_new_block[110]), .D(round_key[110]), .Z(n873[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam xor_56_i4_2_lut_4_lut.init = 16'h6996;
    LUT4 new_block_127__I_0_i113_2_lut (.A(dec_new_block[112]), .B(round_key[112]), 
         .Z(block_new_127__N_1901[112])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i113_2_lut.init = 16'h6666;
    LUT4 i2_2_lut_3_lut_4_lut_adj_217 (.A(block_new_127__N_1901[101]), .B(n33839), 
         .C(n33838), .D(n33837), .Z(n7_adj_7788)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i2_2_lut_3_lut_4_lut_adj_217.init = 16'h6996;
    LUT4 i1_2_lut_rep_405_3_lut (.A(block_new_127__N_1901[58]), .B(block_new_127__N_1901[63]), 
         .C(block_new_127__N_1901[51]), .Z(n33709)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_405_3_lut.init = 16'h9696;
    LUT4 xor_31_i4_2_lut_4_lut (.A(dec_new_block[121]), .B(round_key[121]), 
         .C(dec_new_block[126]), .D(round_key[126]), .Z(n648[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam xor_31_i4_2_lut_4_lut.init = 16'h6996;
    LUT4 xor_636_i4_2_lut_rep_511_4_lut (.A(dec_new_block[17]), .B(round_key[17]), 
         .C(dec_new_block[22]), .D(round_key[22]), .Z(n33815)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam xor_636_i4_2_lut_rep_511_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_4_lut_adj_218 (.A(dec_new_block[110]), .B(round_key[110]), 
         .C(dec_new_block[126]), .D(round_key[126]), .Z(n29339)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_4_lut_adj_218.init = 16'h6996;
    LUT4 i1_4_lut_adj_219 (.A(dec_ctrl_new_2__N_2032), .B(n33842), .C(n20708), 
         .D(n33844), .Z(block_w0_we)) /* synthesis lut_function=(!(A+!(B (C+(D))+!B !((D)+!C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(462[7] 518[14])
    defparam i1_4_lut_adj_219.init = 16'h4450;
    LUT4 block_127__I_0_i48_2_lut (.A(\block_reg[2] [15]), .B(round_key[47]), 
         .Z(block_new_127__N_1645_c[47])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i48_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i47_2_lut (.A(\block_reg[2] [14]), .B(round_key[46]), 
         .Z(block_new_127__N_1645_c[46])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i47_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i111_2_lut (.A(dec_new_block[110]), .B(round_key[110]), 
         .Z(block_new_127__N_1901[110])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i111_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i46_2_lut (.A(\block_reg[2] [13]), .B(round_key[45]), 
         .Z(block_new_127__N_1645_c[45])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i46_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i110_2_lut (.A(dec_new_block[109]), .B(round_key[109]), 
         .Z(block_new_127__N_1901[109])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i110_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i45_2_lut (.A(\block_reg[2] [12]), .B(round_key[44]), 
         .Z(\block_new_127__N_1645[44] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i45_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i44_2_lut (.A(\block_reg[2] [11]), .B(round_key[43]), 
         .Z(\block_new_127__N_1645[43] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i44_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i108_2_lut (.A(dec_new_block[107]), .B(round_key[107]), 
         .Z(block_new_127__N_1901[107])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i108_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i43_2_lut (.A(\block_reg[2] [10]), .B(round_key[42]), 
         .Z(block_new_127__N_1645_c[42])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i43_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i107_2_lut (.A(dec_new_block[106]), .B(round_key[106]), 
         .Z(block_new_127__N_1901[106])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i107_2_lut.init = 16'h6666;
    LUT4 xor_509_i4_2_lut_rep_510_4_lut (.A(dec_new_block[42]), .B(round_key[42]), 
         .C(dec_new_block[47]), .D(round_key[47]), .Z(n33814)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam xor_509_i4_2_lut_rep_510_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_509_4_lut (.A(dec_new_block[39]), .B(round_key[39]), 
         .C(dec_new_block[40]), .D(round_key[40]), .Z(n33813)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_509_4_lut.init = 16'h6996;
    LUT4 new_block_127__I_0_i103_2_lut (.A(dec_new_block[102]), .B(round_key[102]), 
         .Z(block_new_127__N_1901[102])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i103_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i42_2_lut (.A(\block_reg[2] [9]), .B(round_key[41]), 
         .Z(\block_new_127__N_1645[41] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i42_2_lut.init = 16'h6666;
    LUT4 i1_2_lut_rep_508_4_lut (.A(dec_new_block[45]), .B(round_key[45]), 
         .C(dec_new_block[61]), .D(round_key[61]), .Z(n33812)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_rep_508_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_3_lut_adj_220 (.A(block_new_127__N_1901[50]), .B(block_new_127__N_1901[55]), 
         .C(block_new_127__N_1901[43]), .Z(n5_adj_7965)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_3_lut_adj_220.init = 16'h9696;
    LUT4 i1_2_lut_rep_507_4_lut (.A(dec_new_block[37]), .B(round_key[37]), 
         .C(dec_new_block[32]), .D(round_key[32]), .Z(n33811)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_507_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_506_4_lut (.A(dec_new_block[63]), .B(round_key[63]), 
         .C(dec_new_block[56]), .D(round_key[56]), .Z(n33810)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_506_4_lut.init = 16'h6996;
    LUT4 i24_3_lut_4_lut_4_lut (.A(dec_round_nr_c[1]), .B(dec_round_nr[0]), 
         .C(dec_round_nr_c[2]), .D(dec_ctrl_new_2__N_2032), .Z(n14919)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B (C+(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(99[18:30])
    defparam i24_3_lut_4_lut_4_lut.init = 16'h00e1;
    LUT4 i27_3_lut_4_lut_4_lut (.A(dec_round_nr_c[1]), .B(dec_round_nr[0]), 
         .C(dec_round_nr_c[2]), .D(dec_ctrl_new_2__N_2032), .Z(n14930)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B ((D)+!C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(99[18:30])
    defparam i27_3_lut_4_lut_4_lut.init = 16'hffe1;
    LUT4 xor_351_i4_2_lut_rep_505_4_lut (.A(dec_new_block[90]), .B(round_key[90]), 
         .C(dec_new_block[95]), .D(round_key[95]), .Z(n33809)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam xor_351_i4_2_lut_rep_505_4_lut.init = 16'h6996;
    LUT4 i3_3_lut_4_lut_adj_221 (.A(n11890), .B(n29408), .C(n5085[3]), 
         .D(block_new_127__N_1901[51]), .Z(n8_adj_7976)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i3_3_lut_4_lut_adj_221.init = 16'h6996;
    LUT4 xor_43_i5_2_lut_rep_504_4_lut (.A(dec_new_block[115]), .B(round_key[115]), 
         .C(dec_new_block[119]), .D(round_key[119]), .Z(n33808)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam xor_43_i5_2_lut_rep_504_4_lut.init = 16'h6996;
    LUT4 xor_67_i5_2_lut_rep_503_4_lut (.A(dec_new_block[99]), .B(round_key[99]), 
         .C(dec_new_block[103]), .D(round_key[103]), .Z(n33807)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam xor_67_i5_2_lut_rep_503_4_lut.init = 16'h6996;
    LUT4 xor_501_i4_2_lut_rep_502_4_lut (.A(dec_new_block[50]), .B(round_key[50]), 
         .C(dec_new_block[55]), .D(round_key[55]), .Z(n33806)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam xor_501_i4_2_lut_rep_502_4_lut.init = 16'h6996;
    LUT4 xor_489_i4_2_lut_rep_501_4_lut (.A(dec_new_block[58]), .B(round_key[58]), 
         .C(dec_new_block[63]), .D(round_key[63]), .Z(n33805)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam xor_489_i4_2_lut_rep_501_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_500_4_lut (.A(dec_new_block[69]), .B(round_key[69]), 
         .C(dec_new_block[85]), .D(round_key[85]), .Z(n33804)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_500_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_499_4_lut (.A(dec_new_block[93]), .B(round_key[93]), 
         .C(dec_new_block[77]), .D(round_key[77]), .Z(n33803)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_rep_499_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_498_4_lut (.A(dec_new_block[53]), .B(round_key[53]), 
         .C(dec_new_block[61]), .D(round_key[61]), .Z(n33802)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_rep_498_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_497_4_lut (.A(dec_new_block[62]), .B(round_key[62]), 
         .C(dec_new_block[46]), .D(round_key[46]), .Z(n33801)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_rep_497_4_lut.init = 16'h6996;
    LUT4 n2755_bdd_4_lut (.A(n2752[29]), .B(n9422), .C(n30146), .D(n25333), 
         .Z(tmp_sboxw[29])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n2755_bdd_4_lut.init = 16'h00ca;
    LUT4 i1_2_lut_rep_496_4_lut (.A(dec_new_block[60]), .B(round_key[60]), 
         .C(dec_new_block[52]), .D(round_key[52]), .Z(n33800)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_rep_496_4_lut.init = 16'h6996;
    FD1P3AX dec_ctrl_reg_FSM_i0_i1 (.D(n2886), .SP(dec_ctrl_we), .CK(clk_c), 
            .Q(n6363[1]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(462[7] 518[14])
    defparam dec_ctrl_reg_FSM_i0_i1.GSR = "ENABLED";
    LUT4 xor_524_i5_2_lut_rep_495_4_lut (.A(dec_new_block[35]), .B(round_key[35]), 
         .C(dec_new_block[39]), .D(round_key[39]), .Z(n33799)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam xor_524_i5_2_lut_rep_495_4_lut.init = 16'h6996;
    LUT4 xor_509_i5_2_lut_rep_494_4_lut (.A(dec_new_block[43]), .B(round_key[43]), 
         .C(dec_new_block[47]), .D(round_key[47]), .Z(n33798)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam xor_509_i5_2_lut_rep_494_4_lut.init = 16'h6996;
    LUT4 xor_382_i5_2_lut_rep_493_4_lut (.A(dec_new_block[67]), .B(round_key[67]), 
         .C(dec_new_block[71]), .D(round_key[71]), .Z(n33797)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam xor_382_i5_2_lut_rep_493_4_lut.init = 16'h6996;
    LUT4 i2_2_lut_rep_492_4_lut (.A(dec_new_block[70]), .B(round_key[70]), 
         .C(dec_new_block[86]), .D(round_key[86]), .Z(n33796)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i2_2_lut_rep_492_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_491_4_lut (.A(dec_new_block[78]), .B(round_key[78]), 
         .C(dec_new_block[94]), .D(round_key[94]), .Z(n33795)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_rep_491_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_490_4_lut (.A(dec_new_block[84]), .B(round_key[84]), 
         .C(dec_new_block[92]), .D(round_key[92]), .Z(n33794)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_rep_490_4_lut.init = 16'h6996;
    LUT4 xor_351_i5_2_lut_rep_489_4_lut (.A(dec_new_block[91]), .B(round_key[91]), 
         .C(dec_new_block[95]), .D(round_key[95]), .Z(n33793)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam xor_351_i5_2_lut_rep_489_4_lut.init = 16'h6996;
    LUT4 xor_374_i5_2_lut_rep_488_4_lut (.A(dec_new_block[75]), .B(round_key[75]), 
         .C(dec_new_block[79]), .D(round_key[79]), .Z(n33792)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam xor_374_i5_2_lut_rep_488_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_486_4_lut (.A(dec_new_block[118]), .B(round_key[118]), 
         .C(dec_new_block[108]), .D(round_key[108]), .Z(n33790)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_rep_486_4_lut.init = 16'h6996;
    LUT4 xor_649_i5_2_lut_rep_485_4_lut (.A(dec_new_block[11]), .B(round_key[11]), 
         .C(dec_new_block[15]), .D(round_key[15]), .Z(n33789)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam xor_649_i5_2_lut_rep_485_4_lut.init = 16'h6996;
    LUT4 xor_660_i5_2_lut_rep_484_4_lut (.A(dec_new_block[3]), .B(round_key[3]), 
         .C(dec_new_block[7]), .D(round_key[7]), .Z(n33788)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam xor_660_i5_2_lut_rep_484_4_lut.init = 16'h6996;
    LUT4 xor_501_i5_2_lut_rep_483_4_lut (.A(dec_new_block[51]), .B(round_key[51]), 
         .C(dec_new_block[55]), .D(round_key[55]), .Z(n33787)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam xor_501_i5_2_lut_rep_483_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_482_4_lut (.A(dec_new_block[38]), .B(round_key[38]), 
         .C(dec_new_block[54]), .D(round_key[54]), .Z(n33786)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_482_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_481_4_lut (.A(dec_new_block[76]), .B(round_key[76]), 
         .C(dec_new_block[68]), .D(round_key[68]), .Z(n33785)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_rep_481_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_480_4_lut (.A(dec_new_block[22]), .B(round_key[22]), 
         .C(dec_new_block[6]), .D(round_key[6]), .Z(n33784)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_rep_480_4_lut.init = 16'h6996;
    LUT4 xor_627_i5_2_lut_rep_479_4_lut (.A(dec_new_block[27]), .B(round_key[27]), 
         .C(dec_new_block[31]), .D(round_key[31]), .Z(n33783)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam xor_627_i5_2_lut_rep_479_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_478_4_lut (.A(dec_new_block[20]), .B(round_key[20]), 
         .C(dec_new_block[12]), .D(round_key[12]), .Z(n33782)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_rep_478_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_477_4_lut (.A(dec_new_block[17]), .B(round_key[17]), 
         .C(dec_new_block[9]), .D(round_key[9]), .Z(n33781)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_rep_477_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_476_4_lut (.A(dec_new_block[29]), .B(round_key[29]), 
         .C(dec_new_block[13]), .D(round_key[13]), .Z(n33780)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_476_4_lut.init = 16'h6996;
    LUT4 n2756_bdd_4_lut (.A(n2752[28]), .B(n9420), .C(n30146), .D(n25333), 
         .Z(tmp_sboxw[28])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n2756_bdd_4_lut.init = 16'h00ca;
    LUT4 i1_2_lut_rep_475_4_lut (.A(dec_new_block[5]), .B(round_key[5]), 
         .C(dec_new_block[21]), .D(round_key[21]), .Z(n33779)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_rep_475_4_lut.init = 16'h6996;
    LUT4 i3_3_lut_4_lut_adj_222 (.A(block_new_127__N_1901[48]), .B(n33670), 
         .C(n33812), .D(block_new_127__N_1901[55]), .Z(n8_adj_7728)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i3_3_lut_4_lut_adj_222.init = 16'h6996;
    LUT4 xor_634_i5_2_lut_rep_474_4_lut (.A(dec_new_block[19]), .B(round_key[19]), 
         .C(dec_new_block[23]), .D(round_key[23]), .Z(n33778)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam xor_634_i5_2_lut_rep_474_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_473_4_lut (.A(dec_new_block[25]), .B(round_key[25]), 
         .C(dec_new_block[17]), .D(round_key[17]), .Z(n33777)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_473_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_471_4_lut (.A(dec_new_block[23]), .B(round_key[23]), 
         .C(dec_new_block[24]), .D(round_key[24]), .Z(n33775)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_rep_471_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_470_4_lut (.A(dec_new_block[14]), .B(round_key[14]), 
         .C(dec_new_block[22]), .D(round_key[22]), .Z(n33774)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_470_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_469_4_lut (.A(dec_new_block[31]), .B(round_key[31]), 
         .C(dec_new_block[8]), .D(round_key[8]), .Z(n33773)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_rep_469_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_468_4_lut (.A(dec_new_block[47]), .B(round_key[47]), 
         .C(dec_new_block[56]), .D(round_key[56]), .Z(n33772)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_468_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_467_4_lut (.A(dec_new_block[64]), .B(round_key[64]), 
         .C(dec_new_block[80]), .D(round_key[80]), .Z(n33771)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_rep_467_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_466_4_lut (.A(dec_new_block[109]), .B(round_key[109]), 
         .C(dec_new_block[108]), .D(round_key[108]), .Z(n33770)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_rep_466_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_465_4_lut (.A(dec_new_block[110]), .B(round_key[110]), 
         .C(dec_new_block[102]), .D(round_key[102]), .Z(n33769)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_rep_465_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_464_4_lut (.A(dec_new_block[103]), .B(round_key[103]), 
         .C(dec_new_block[104]), .D(round_key[104]), .Z(n33768)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_rep_464_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_463_4_lut (.A(dec_new_block[119]), .B(round_key[119]), 
         .C(dec_new_block[120]), .D(round_key[120]), .Z(n33767)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_463_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_462_4_lut (.A(dec_new_block[102]), .B(round_key[102]), 
         .C(dec_new_block[118]), .D(round_key[118]), .Z(n33766)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_462_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_461_4_lut (.A(dec_new_block[9]), .B(round_key[9]), 
         .C(dec_new_block[1]), .D(round_key[1]), .Z(n33765)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_461_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_460_4_lut (.A(dec_new_block[46]), .B(round_key[46]), 
         .C(dec_new_block[55]), .D(round_key[55]), .Z(n33764)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_460_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_459_4_lut (.A(dec_new_block[44]), .B(round_key[44]), 
         .C(dec_new_block[36]), .D(round_key[36]), .Z(n33763)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_rep_459_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_458_4_lut (.A(dec_new_block[86]), .B(round_key[86]), 
         .C(dec_new_block[78]), .D(round_key[78]), .Z(n33762)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_458_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_457_4_lut (.A(dec_new_block[5]), .B(round_key[5]), 
         .C(dec_new_block[4]), .D(round_key[4]), .Z(n33761)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_rep_457_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_456_4_lut (.A(dec_new_block[47]), .B(round_key[47]), 
         .C(dec_new_block[46]), .D(round_key[46]), .Z(n33760)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_rep_456_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_455_4_lut (.A(dec_new_block[98]), .B(round_key[98]), 
         .C(dec_new_block[122]), .D(round_key[122]), .Z(n33759)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_455_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_454_4_lut (.A(dec_new_block[121]), .B(round_key[121]), 
         .C(dec_new_block[96]), .D(round_key[96]), .Z(n33758)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_454_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_453_4_lut (.A(dec_new_block[30]), .B(round_key[30]), 
         .C(dec_new_block[15]), .D(round_key[15]), .Z(n33757)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_rep_453_4_lut.init = 16'h6996;
    FD1P3AX sword_ctr_reg_FSM_i0_i3 (.D(n2689[3]), .SP(sword_ctr_we), .CK(clk_c), 
            .Q(n6362[3]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam sword_ctr_reg_FSM_i0_i3.GSR = "ENABLED";
    FD1P3AX sword_ctr_reg_FSM_i0_i2 (.D(n2689[2]), .SP(sword_ctr_we), .CK(clk_c), 
            .Q(n6362[2]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam sword_ctr_reg_FSM_i0_i2.GSR = "ENABLED";
    FD1P3IX sword_ctr_reg_FSM_i0_i1 (.D(n6362[0]), .SP(sword_ctr_we), .CD(n33909), 
            .CK(clk_c), .Q(n6362[1]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam sword_ctr_reg_FSM_i0_i1.GSR = "ENABLED";
    FD1P3AX dec_ctrl_reg_FSM_i0_i2 (.D(n33858), .SP(dec_ctrl_we), .CK(clk_c), 
            .Q(n6363[2]));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(462[7] 518[14])
    defparam dec_ctrl_reg_FSM_i0_i2.GSR = "ENABLED";
    FD1P3AY dec_ctrl_reg_FSM_i0_i3 (.D(n28836), .SP(dec_ctrl_we), .CK(clk_c), 
            .Q(dec_ctrl_new_2__N_2032));   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(462[7] 518[14])
    defparam dec_ctrl_reg_FSM_i0_i3.GSR = "ENABLED";
    PFUMX mux_625_i126 (.BLUT(n2_adj_7997), .ALUT(n4540[125]), .C0(n30026), 
          .Z(n3899[125]));
    PFUMX mux_625_i124 (.BLUT(n2_adj_7995), .ALUT(n4540[123]), .C0(n30026), 
          .Z(n3899[123]));
    PFUMX mux_625_i84 (.BLUT(n2_adj_7993), .ALUT(n4540[83]), .C0(n30026), 
          .Z(n3899[83]));
    PFUMX mux_625_i76 (.BLUT(n2_adj_7991), .ALUT(n4540[75]), .C0(n30026), 
          .Z(n3899[75]));
    LUT4 i1_2_lut_rep_545_4_lut (.A(dec_round_nr_c[3]), .B(n33936), .C(dec_round_nr_c[2]), 
         .D(n6363[1]), .Z(n33849)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_545_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_4_lut_adj_223 (.A(dec_round_nr_c[3]), .B(n33936), .C(dec_round_nr_c[2]), 
         .D(n6363[0]), .Z(n14890)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_2_lut_4_lut_adj_223.init = 16'h0100;
    PFUMX mux_625_i52 (.BLUT(n2_adj_7989), .ALUT(n4540[51]), .C0(n30026), 
          .Z(n3899[51]));
    PFUMX mux_625_i28 (.BLUT(n2_adj_7986), .ALUT(n4540[27]), .C0(n30026), 
          .Z(n3899[27]));
    PFUMX mux_625_i12 (.BLUT(n2_adj_7983), .ALUT(n4540[11]), .C0(n30026), 
          .Z(n3899[11]));
    PFUMX mux_625_i116 (.BLUT(n2_adj_7980), .ALUT(n4540[115]), .C0(n30026), 
          .Z(n3899[115]));
    PFUMX mux_625_i108 (.BLUT(n2_adj_7977), .ALUT(n4540[107]), .C0(n30026), 
          .Z(n3899[107]));
    PFUMX mux_625_i106 (.BLUT(n2_adj_7974), .ALUT(n4540[105]), .C0(n30026), 
          .Z(n3899[105]));
    PFUMX mux_625_i92 (.BLUT(n2_adj_7972), .ALUT(n4540[91]), .C0(n30026), 
          .Z(n3899[91]));
    PFUMX mux_625_i86 (.BLUT(n2_adj_7970), .ALUT(n4540[85]), .C0(n30026), 
          .Z(n3899[85]));
    PFUMX mux_625_i60 (.BLUT(n2_adj_7967), .ALUT(n4540[59]), .C0(n30026), 
          .Z(n3899[59]));
    PFUMX mux_625_i50 (.BLUT(n2_adj_7964), .ALUT(n4540[49]), .C0(n30026), 
          .Z(n3899[49]));
    PFUMX mux_625_i44 (.BLUT(n2_adj_7962), .ALUT(n4540[43]), .C0(n30026), 
          .Z(n3899[43]));
    PFUMX mux_625_i6 (.BLUT(n2_adj_7960), .ALUT(n4540[5]), .C0(n30026), 
          .Z(n3899[5]));
    PFUMX mux_625_i109 (.BLUT(n2_adj_7957), .ALUT(n4540[108]), .C0(n30026), 
          .Z(n3899[108]));
    PFUMX mux_625_i102 (.BLUT(n2_adj_7954), .ALUT(n4540[101]), .C0(n30026), 
          .Z(n3899[101]));
    PFUMX mux_625_i101 (.BLUT(n2_adj_7951), .ALUT(n4540[100]), .C0(n30026), 
          .Z(n3899[100]));
    PFUMX mux_625_i100 (.BLUT(n2_adj_7948), .ALUT(n4540[99]), .C0(n30026), 
          .Z(n3899[99]));
    PFUMX mux_625_i94 (.BLUT(n2_adj_7945), .ALUT(n4540[93]), .C0(n30026), 
          .Z(n3899[93]));
    PFUMX mux_625_i93 (.BLUT(n2_adj_7942), .ALUT(n4540[92]), .C0(n30026), 
          .Z(n3899[92]));
    PFUMX mux_625_i85 (.BLUT(n2_adj_7940), .ALUT(n4540[84]), .C0(n30026), 
          .Z(n3899[84]));
    PFUMX mux_625_i77 (.BLUT(n2_adj_7938), .ALUT(n4540[76]), .C0(n30026), 
          .Z(n3899[76]));
    PFUMX mux_625_i70 (.BLUT(n2_adj_7935), .ALUT(n4540[69]), .C0(n30026), 
          .Z(n3899[69]));
    PFUMX mux_625_i65 (.BLUT(n2_adj_7933), .ALUT(n4540[64]), .C0(n30026), 
          .Z(n3899[64]));
    PFUMX mux_625_i62 (.BLUT(n2_adj_7931), .ALUT(n4540[61]), .C0(n30026), 
          .Z(n3899[61]));
    PFUMX mux_625_i54 (.BLUT(n2_adj_7930), .ALUT(n4540[53]), .C0(n30026), 
          .Z(n3899[53]));
    PFUMX mux_625_i53 (.BLUT(n2_adj_7928), .ALUT(n4540[52]), .C0(n30026), 
          .Z(n3899[52]));
    PFUMX mux_625_i46 (.BLUT(n2_adj_7925), .ALUT(n4540[45]), .C0(n30026), 
          .Z(n3899[45]));
    PFUMX mux_625_i45 (.BLUT(n2_adj_7922), .ALUT(n4540[44]), .C0(n30026), 
          .Z(n3899[44]));
    PFUMX mux_625_i37 (.BLUT(n2_adj_7920), .ALUT(n4540[36]), .C0(n30026), 
          .Z(n3899[36]));
    PFUMX mux_625_i36 (.BLUT(n2_adj_7917), .ALUT(n4540[35]), .C0(n30026), 
          .Z(n3899[35]));
    PFUMX mux_625_i34 (.BLUT(n2_adj_7914), .ALUT(n4540[33]), .C0(n30026), 
          .Z(n3899[33]));
    PFUMX mux_625_i30 (.BLUT(n2_adj_7912), .ALUT(n4540[29]), .C0(n30026), 
          .Z(n3899[29]));
    PFUMX mux_625_i29 (.BLUT(n2_adj_7910), .ALUT(n4540[28]), .C0(n30026), 
          .Z(n3899[28]));
    PFUMX mux_625_i27 (.BLUT(n2_adj_7906), .ALUT(n4540[26]), .C0(n30026), 
          .Z(n3899[26]));
    PFUMX mux_625_i25 (.BLUT(n2_adj_7904), .ALUT(n4540[24]), .C0(n30026), 
          .Z(n3899[24]));
    PFUMX mux_625_i20 (.BLUT(n2_adj_7903), .ALUT(n4540[19]), .C0(n30026), 
          .Z(n3899[19]));
    PFUMX mux_625_i17 (.BLUT(n2_adj_7900), .ALUT(n4540[16]), .C0(n30026), 
          .Z(n3899[16]));
    PFUMX mux_625_i13 (.BLUT(n2_adj_7898), .ALUT(n4540[12]), .C0(n30026), 
          .Z(n3899[12]));
    PFUMX mux_625_i9 (.BLUT(n2_adj_7894), .ALUT(n4540[8]), .C0(n30026), 
          .Z(n3899[8]));
    PFUMX mux_625_i5 (.BLUT(n2_adj_7892), .ALUT(n4540[4]), .C0(n30026), 
          .Z(n3899[4]));
    PFUMX mux_625_i4 (.BLUT(n2_adj_7890), .ALUT(n4540[3]), .C0(n30026), 
          .Z(n3899[3]));
    PFUMX mux_625_i128 (.BLUT(n2_adj_7887), .ALUT(n4540[127]), .C0(n30026), 
          .Z(n3899[127]));
    PFUMX mux_625_i127 (.BLUT(n2_adj_7884), .ALUT(n4540[126]), .C0(n30026), 
          .Z(n3899[126]));
    PFUMX mux_625_i125 (.BLUT(n2_adj_7882), .ALUT(n4540[124]), .C0(n30026), 
          .Z(n3899[124]));
    PFUMX mux_625_i123 (.BLUT(n2_adj_7879), .ALUT(n4540[122]), .C0(n30026), 
          .Z(n3899[122]));
    PFUMX mux_625_i119 (.BLUT(n2_adj_7876), .ALUT(n4540[118]), .C0(n30026), 
          .Z(n3899[118]));
    PFUMX mux_625_i118 (.BLUT(n2_adj_7873), .ALUT(n4540[117]), .C0(n30026), 
          .Z(n3899[117]));
    PFUMX mux_625_i117 (.BLUT(n2_adj_7870), .ALUT(n4540[116]), .C0(n30026), 
          .Z(n3899[116]));
    PFUMX mux_625_i114 (.BLUT(n2_adj_7868), .ALUT(n4540[113]), .C0(n30026), 
          .Z(n3899[113]));
    PFUMX mux_625_i112 (.BLUT(n2_adj_7865), .ALUT(n4540[111]), .C0(n30026), 
          .Z(n3899[111]));
    PFUMX mux_625_i110 (.BLUT(n2_adj_7863), .ALUT(n4540[109]), .C0(n30026), 
          .Z(n3899[109]));
    PFUMX mux_625_i103 (.BLUT(n2_adj_7861), .ALUT(n4540[102]), .C0(n30026), 
          .Z(n3899[102]));
    PFUMX mux_625_i96 (.BLUT(n2_adj_7859), .ALUT(n4540[95]), .C0(n30026), 
          .Z(n3899[95]));
    PFUMX mux_625_i95 (.BLUT(n2_adj_7857), .ALUT(n4540[94]), .C0(n30026), 
          .Z(n3899[94]));
    PFUMX mux_625_i91 (.BLUT(n2_adj_7855), .ALUT(n4540[90]), .C0(n30026), 
          .Z(n3899[90]));
    PFUMX mux_625_i89 (.BLUT(n2_adj_7852), .ALUT(n4540[88]), .C0(n30026), 
          .Z(n3899[88]));
    PFUMX mux_625_i82 (.BLUT(n2_adj_7849), .ALUT(n4540[81]), .C0(n30026), 
          .Z(n3899[81]));
    PFUMX mux_625_i79 (.BLUT(n2_adj_7846), .ALUT(n4540[78]), .C0(n30026), 
          .Z(n3899[78]));
    PFUMX mux_625_i78 (.BLUT(n2_adj_7842), .ALUT(n4540[77]), .C0(n30026), 
          .Z(n3899[77]));
    PFUMX mux_625_i75 (.BLUT(n2_adj_7840), .ALUT(n4540[74]), .C0(n30026), 
          .Z(n3899[74]));
    PFUMX mux_625_i69 (.BLUT(n2_adj_7838), .ALUT(n4540[68]), .C0(n30026), 
          .Z(n3899[68]));
    PFUMX mux_625_i68 (.BLUT(n2_adj_7835), .ALUT(n4540[67]), .C0(n30026), 
          .Z(n3899[67]));
    PFUMX mux_625_i67 (.BLUT(n2_adj_7832), .ALUT(n4540[66]), .C0(n30026), 
          .Z(n3899[66]));
    PFUMX mux_625_i61 (.BLUT(n2_adj_7828), .ALUT(n4540[60]), .C0(n30026), 
          .Z(n3899[60]));
    PFUMX mux_625_i48 (.BLUT(n2_adj_7827), .ALUT(n4540[47]), .C0(n30026), 
          .Z(n3899[47]));
    PFUMX mux_625_i43 (.BLUT(n2_adj_7825), .ALUT(n4540[42]), .C0(n30026), 
          .Z(n3899[42]));
    PFUMX mux_625_i42 (.BLUT(n2_adj_7823), .ALUT(n4540[41]), .C0(n30026), 
          .Z(n3899[41]));
    PFUMX mux_625_i39 (.BLUT(n2_adj_7819), .ALUT(n4540[38]), .C0(n30026), 
          .Z(n3899[38]));
    PFUMX mux_625_i38 (.BLUT(n2_adj_7815), .ALUT(n4540[37]), .C0(n30026), 
          .Z(n3899[37]));
    PFUMX mux_625_i32 (.BLUT(n2_adj_7811), .ALUT(n4540[31]), .C0(n30026), 
          .Z(n3899[31]));
    PFUMX mux_625_i31 (.BLUT(n2_adj_7808), .ALUT(n4540[30]), .C0(n30026), 
          .Z(n3899[30]));
    PFUMX mux_625_i22 (.BLUT(n2_adj_7805), .ALUT(n4540[21]), .C0(n30026), 
          .Z(n3899[21]));
    PFUMX mux_625_i21 (.BLUT(n2_adj_7801), .ALUT(n4540[20]), .C0(n30026), 
          .Z(n3899[20]));
    PFUMX mux_625_i15 (.BLUT(n2_adj_7798), .ALUT(n4540[14]), .C0(n30026), 
          .Z(n3899[14]));
    PFUMX mux_625_i11 (.BLUT(n2_adj_7796), .ALUT(n4540[10]), .C0(n30026), 
          .Z(n3899[10]));
    PFUMX mux_625_i10 (.BLUT(n2_adj_7793), .ALUT(n4540[9]), .C0(n30026), 
          .Z(n3899[9]));
    PFUMX mux_625_i7 (.BLUT(n2_adj_7790), .ALUT(n4540[6]), .C0(n30026), 
          .Z(n3899[6]));
    PFUMX mux_625_i3 (.BLUT(n2_adj_7787), .ALUT(n4540[2]), .C0(n30026), 
          .Z(n3899[2]));
    PFUMX mux_625_i1 (.BLUT(n2_adj_7784), .ALUT(n4540[0]), .C0(n30026), 
          .Z(n3899[0]));
    PFUMX mux_625_i122 (.BLUT(n2_adj_7783), .ALUT(n4540[121]), .C0(n30026), 
          .Z(n3899[121]));
    PFUMX mux_625_i121 (.BLUT(n2_adj_7781), .ALUT(n4540[120]), .C0(n30026), 
          .Z(n3899[120]));
    PFUMX mux_625_i113 (.BLUT(n2_adj_7779), .ALUT(n4540[112]), .C0(n30026), 
          .Z(n3899[112]));
    PFUMX mux_625_i111 (.BLUT(n2_adj_7776), .ALUT(n4540[110]), .C0(n30026), 
          .Z(n3899[110]));
    PFUMX mux_625_i107 (.BLUT(n2_adj_7773), .ALUT(n4540[106]), .C0(n30026), 
          .Z(n3899[106]));
    PFUMX mux_625_i105 (.BLUT(n2_adj_7772), .ALUT(n4540[104]), .C0(n30026), 
          .Z(n3899[104]));
    PFUMX mux_625_i104 (.BLUT(n2_adj_7770), .ALUT(n4540[103]), .C0(n30026), 
          .Z(n3899[103]));
    PFUMX mux_625_i99 (.BLUT(n2_adj_7767), .ALUT(n4540[98]), .C0(n30026), 
          .Z(n3899[98]));
    PFUMX mux_625_i98 (.BLUT(n2_adj_7765), .ALUT(n4540[97]), .C0(n30026), 
          .Z(n3899[97]));
    PFUMX mux_625_i97 (.BLUT(n2_adj_7763), .ALUT(n4540[96]), .C0(n30026), 
          .Z(n3899[96]));
    PFUMX mux_625_i90 (.BLUT(n2_adj_7760), .ALUT(n4540[89]), .C0(n30026), 
          .Z(n3899[89]));
    PFUMX mux_625_i87 (.BLUT(n2_adj_7757), .ALUT(n4540[86]), .C0(n30026), 
          .Z(n3899[86]));
    PFUMX mux_625_i83 (.BLUT(n2_adj_7755), .ALUT(n4540[82]), .C0(n30026), 
          .Z(n3899[82]));
    PFUMX mux_625_i81 (.BLUT(n2_adj_7751), .ALUT(n4540[80]), .C0(n30026), 
          .Z(n3899[80]));
    PFUMX mux_625_i80 (.BLUT(n2_adj_7749), .ALUT(n4540[79]), .C0(n30026), 
          .Z(n3899[79]));
    PFUMX mux_625_i74 (.BLUT(n2_adj_7747), .ALUT(n4540[73]), .C0(n30026), 
          .Z(n3899[73]));
    PFUMX mux_625_i72 (.BLUT(n2_adj_7744), .ALUT(n4540[71]), .C0(n30026), 
          .Z(n3899[71]));
    PFUMX mux_625_i71 (.BLUT(n2_adj_7741), .ALUT(n4540[70]), .C0(n30026), 
          .Z(n3899[70]));
    PFUMX mux_625_i64 (.BLUT(n2_adj_7739), .ALUT(n4540[63]), .C0(n30026), 
          .Z(n3899[63]));
    PFUMX mux_625_i63 (.BLUT(n2_adj_7737), .ALUT(n4540[62]), .C0(n30026), 
          .Z(n3899[62]));
    PFUMX mux_625_i58 (.BLUT(n2_adj_7734), .ALUT(n4540[57]), .C0(n30026), 
          .Z(n3899[57]));
    LUT4 new_block_127__I_0_i106_2_lut (.A(dec_new_block[105]), .B(round_key[105]), 
         .Z(block_new_127__N_1901[105])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i106_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i41_2_lut (.A(\block_reg[2] [8]), .B(round_key[40]), 
         .Z(block_new_127__N_1645_c[40])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i41_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i105_2_lut (.A(dec_new_block[104]), .B(round_key[104]), 
         .Z(block_new_127__N_1901[104])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i105_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i72_2_lut (.A(\block_reg[1] [7]), .B(round_key[71]), 
         .Z(\block_new_127__N_1645[71] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i72_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i104_2_lut (.A(dec_new_block[103]), .B(round_key[103]), 
         .Z(block_new_127__N_1901[103])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i104_2_lut.init = 16'h6666;
    PFUMX mux_625_i57 (.BLUT(n2_adj_7729), .ALUT(n4540[56]), .C0(n30026), 
          .Z(n3899[56]));
    PFUMX mux_625_i55 (.BLUT(n2_adj_7726), .ALUT(n4540[54]), .C0(n30026), 
          .Z(n3899[54]));
    PFUMX mux_625_i51 (.BLUT(n2_adj_7723), .ALUT(n4540[50]), .C0(n30026), 
          .Z(n3899[50]));
    PFUMX mux_625_i47 (.BLUT(n2_adj_7721), .ALUT(n4540[46]), .C0(n30026), 
          .Z(n3899[46]));
    LUT4 i29_4_lut_4_lut (.A(n14912), .B(n33942), .C(n149), .D(encdec_reg), 
         .Z(n14933)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(72[15:32])
    defparam i29_4_lut_4_lut.init = 16'ha0ac;
    PFUMX mux_625_i41 (.BLUT(n2_adj_7717), .ALUT(n4540[40]), .C0(n30026), 
          .Z(n3899[40]));
    PFUMX mux_625_i40 (.BLUT(n2_adj_7715), .ALUT(n4540[39]), .C0(n30026), 
          .Z(n3899[39]));
    LUT4 i1_2_lut_rep_605 (.A(n6363[0]), .B(n6363[2]), .Z(n33909)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(462[7] 518[14])
    defparam i1_2_lut_rep_605.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_adj_224 (.A(n6363[0]), .B(n6363[2]), .C(n6363[1]), 
         .Z(sword_ctr_we)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(462[7] 518[14])
    defparam i1_2_lut_3_lut_adj_224.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut_4_lut_adj_225 (.A(block_new_127__N_1901[107]), .B(block_new_127__N_1901[111]), 
         .C(n33714), .D(n33839), .Z(n4_adj_7921)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_3_lut_4_lut_adj_225.init = 16'h6996;
    LUT4 i1_2_lut_3_lut_4_lut_adj_226 (.A(n6363[0]), .B(n6363[2]), .C(n6362[3]), 
         .D(n6363[1]), .Z(n2689[0])) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(462[7] 518[14])
    defparam i1_2_lut_3_lut_4_lut_adj_226.init = 16'hfeff;
    LUT4 i15221_2_lut_3_lut_4_lut (.A(n6363[0]), .B(n6363[2]), .C(n6362[1]), 
         .D(n6363[1]), .Z(n2689[2])) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(462[7] 518[14])
    defparam i15221_2_lut_3_lut_4_lut.init = 16'h1000;
    PFUMX mux_625_i35 (.BLUT(n2_adj_7712), .ALUT(n4540[34]), .C0(n30026), 
          .Z(n3899[34]));
    LUT4 i15222_2_lut_3_lut_4_lut (.A(n6363[0]), .B(n6363[2]), .C(n6362[2]), 
         .D(n6363[1]), .Z(n2689[3])) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(462[7] 518[14])
    defparam i15222_2_lut_3_lut_4_lut.init = 16'h1000;
    PFUMX mux_625_i33 (.BLUT(n2_adj_7710), .ALUT(n4540[32]), .C0(n30026), 
          .Z(n3899[32]));
    PFUMX mux_625_i26 (.BLUT(n2_adj_7708), .ALUT(n4540[25]), .C0(n30026), 
          .Z(n3899[25]));
    PFUMX mux_625_i23 (.BLUT(n2_adj_7706), .ALUT(n4540[22]), .C0(n30026), 
          .Z(n3899[22]));
    LUT4 i1_2_lut_rep_397_3_lut (.A(block_new_127__N_1901[107]), .B(block_new_127__N_1901[111]), 
         .C(block_new_127__N_1901[100]), .Z(n33701)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_397_3_lut.init = 16'h9696;
    PFUMX mux_625_i19 (.BLUT(n2_adj_7705), .ALUT(n4540[18]), .C0(n30026), 
          .Z(n3899[18]));
    LUT4 i1_2_lut_rep_386_3_lut_4_lut (.A(block_new_127__N_1901[107]), .B(block_new_127__N_1901[111]), 
         .C(block_new_127__N_1901[127]), .D(block_new_127__N_1901[123]), 
         .Z(n33690)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_386_3_lut_4_lut.init = 16'h6996;
    LUT4 new_block_127__I_0_i101_2_lut (.A(dec_new_block[100]), .B(round_key[100]), 
         .Z(block_new_127__N_1901[100])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i101_2_lut.init = 16'h6666;
    PFUMX mux_625_i18 (.BLUT(n2_adj_7704), .ALUT(n4540[17]), .C0(n30026), 
          .Z(n3899[17]));
    LUT4 block_127__I_0_i68_2_lut (.A(\block_reg[1] [3]), .B(round_key[67]), 
         .Z(\block_new_127__N_1645[67] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i68_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i100_2_lut (.A(dec_new_block[99]), .B(round_key[99]), 
         .Z(block_new_127__N_1901[99])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i100_2_lut.init = 16'h6666;
    PFUMX mux_625_i16 (.BLUT(n2_adj_7702), .ALUT(n4540[15]), .C0(n30026), 
          .Z(n3899[15]));
    LUT4 block_127__I_0_i67_2_lut (.A(\block_reg[1] [2]), .B(round_key[66]), 
         .Z(block_new_127__N_1645_c[66])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i67_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i99_2_lut (.A(dec_new_block[98]), .B(round_key[98]), 
         .Z(block_new_127__N_1901[98])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i99_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i66_2_lut (.A(\block_reg[1] [1]), .B(round_key[65]), 
         .Z(\block_new_127__N_1645[65] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i66_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i98_2_lut (.A(dec_new_block[97]), .B(round_key[97]), 
         .Z(block_new_127__N_1901[97])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i98_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i65_2_lut (.A(\block_reg[1] [0]), .B(round_key[64]), 
         .Z(\block_new_127__N_1645[64] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i65_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i97_2_lut (.A(dec_new_block[96]), .B(round_key[96]), 
         .Z(block_new_127__N_1901[96])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i97_2_lut.init = 16'h6666;
    PFUMX mux_625_i14 (.BLUT(n2_adj_7698), .ALUT(n4540[13]), .C0(n30026), 
          .Z(n3899[13]));
    LUT4 block_127__I_0_i96_2_lut (.A(\block_reg[1] [31]), .B(round_key[95]), 
         .Z(block_new_127__N_1645_c[95])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i96_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i96_2_lut (.A(dec_new_block[95]), .B(round_key[95]), 
         .Z(block_new_127__N_1901[95])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i96_2_lut.init = 16'h6666;
    PFUMX mux_625_i2 (.BLUT(n2), .ALUT(n4540[1]), .C0(n30026), .Z(n3899[1]));
    LUT4 block_127__I_0_i95_2_lut (.A(\block_reg[1] [30]), .B(round_key[94]), 
         .Z(block_new_127__N_1645_c[94])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i95_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i95_2_lut (.A(dec_new_block[94]), .B(round_key[94]), 
         .Z(block_new_127__N_1901[94])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i95_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i94_2_lut (.A(\block_reg[1] [29]), .B(round_key[93]), 
         .Z(block_new_127__N_1645_c[93])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i94_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i94_2_lut (.A(dec_new_block[93]), .B(round_key[93]), 
         .Z(block_new_127__N_1901[93])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i94_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i93_2_lut (.A(\block_reg[1] [28]), .B(round_key[92]), 
         .Z(\block_new_127__N_1645[92] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i93_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i93_2_lut (.A(dec_new_block[92]), .B(round_key[92]), 
         .Z(block_new_127__N_1901[92])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i93_2_lut.init = 16'h6666;
    LUT4 i27579_3_lut_4_lut (.A(block_new_127__N_1645_c[96]), .B(update_type[0]), 
         .C(n33844), .D(n12933), .Z(n4540[0])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam i27579_3_lut_4_lut.init = 16'hf808;
    LUT4 i2_2_lut_3_lut_4_lut_adj_227 (.A(block_new_127__N_1901[126]), .B(block_new_127__N_1901[111]), 
         .C(n33791), .D(block_new_127__N_1901[109]), .Z(n7_adj_7847)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i2_2_lut_3_lut_4_lut_adj_227.init = 16'h6996;
    LUT4 i2_2_lut_3_lut_adj_228 (.A(block_new_127__N_1901[126]), .B(block_new_127__N_1901[111]), 
         .C(n29231), .Z(n6_adj_7886)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i2_2_lut_3_lut_adj_228.init = 16'h9696;
    LUT4 block_127__I_0_i92_2_lut (.A(\block_reg[1] [27]), .B(round_key[91]), 
         .Z(\block_new_127__N_1645[91] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i92_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i92_2_lut (.A(dec_new_block[91]), .B(round_key[91]), 
         .Z(block_new_127__N_1901[91])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i92_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i91_2_lut (.A(\block_reg[1] [26]), .B(round_key[90]), 
         .Z(block_new_127__N_1645_c[90])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i91_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i91_2_lut (.A(dec_new_block[90]), .B(round_key[90]), 
         .Z(block_new_127__N_1901[90])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i91_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i90_2_lut (.A(\block_reg[1] [25]), .B(round_key[89]), 
         .Z(\block_new_127__N_1645[89] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i90_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i90_2_lut (.A(dec_new_block[89]), .B(round_key[89]), 
         .Z(block_new_127__N_1901[89])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i90_2_lut.init = 16'h6666;
    LUT4 i1_2_lut_rep_631 (.A(dec_ctrl_new_2__N_2032), .B(n6363[2]), .Z(n33935)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_631.init = 16'heeee;
    LUT4 i27866_2_lut_2_lut_3_lut_3_lut_2_lut_3_lut_4_lut (.A(dec_ctrl_new_2__N_2032), 
         .B(n6363[2]), .C(n33856), .D(n6363[1]), .Z(n30026)) /* synthesis lut_function=(A+(B+!(C+(D)))) */ ;
    defparam i27866_2_lut_2_lut_3_lut_3_lut_2_lut_3_lut_4_lut.init = 16'heeef;
    LUT4 i2_2_lut_3_lut_adj_229 (.A(block_new_127__N_1901[57]), .B(block_new_127__N_1901[49]), 
         .C(block_new_127__N_1901[33]), .Z(n7_adj_7973)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i2_2_lut_3_lut_adj_229.init = 16'h9696;
    LUT4 block_127__I_0_i89_2_lut (.A(\block_reg[1] [24]), .B(round_key[88]), 
         .Z(block_new_127__N_1645_c[88])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i89_2_lut.init = 16'h6666;
    LUT4 i27882_2_lut_rep_540_2_lut_3_lut_4_lut (.A(dec_ctrl_new_2__N_2032), 
         .B(n6363[2]), .C(n33856), .D(n6363[1]), .Z(n33844)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i27882_2_lut_rep_540_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 new_block_127__I_0_i89_2_lut (.A(dec_new_block[88]), .B(round_key[88]), 
         .Z(block_new_127__N_1901[88])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i89_2_lut.init = 16'h6666;
    LUT4 i15231_2_lut_rep_632 (.A(dec_round_nr_c[1]), .B(dec_round_nr[0]), 
         .Z(n33936)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(99[18:30])
    defparam i15231_2_lut_rep_632.init = 16'heeee;
    LUT4 i2_3_lut_rep_552_4_lut (.A(dec_round_nr_c[1]), .B(dec_round_nr[0]), 
         .C(dec_round_nr_c[2]), .D(dec_round_nr_c[3]), .Z(n33856)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(99[18:30])
    defparam i2_3_lut_rep_552_4_lut.init = 16'hfffe;
    LUT4 block_127__I_0_i120_2_lut (.A(\block_reg[0] [23]), .B(round_key[119]), 
         .Z(\block_new_127__N_1645[119] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i120_2_lut.init = 16'h6666;
    LUT4 i15232_3_lut_4_lut (.A(dec_round_nr_c[1]), .B(dec_round_nr[0]), 
         .C(dec_round_nr_c[3]), .D(dec_round_nr_c[2]), .Z(n14939)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)+!C !(D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_core.v(99[18:30])
    defparam i15232_3_lut_4_lut.init = 16'hf0e1;
    LUT4 new_block_127__I_0_i88_2_lut (.A(dec_new_block[87]), .B(round_key[87]), 
         .Z(block_new_127__N_1901[87])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i88_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i119_2_lut (.A(\block_reg[0] [22]), .B(round_key[118]), 
         .Z(\block_new_127__N_1645[118] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i119_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i87_2_lut (.A(dec_new_block[86]), .B(round_key[86]), 
         .Z(block_new_127__N_1901[86])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i87_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i118_2_lut (.A(\block_reg[0] [21]), .B(round_key[117]), 
         .Z(block_new_127__N_1645_c[117])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i118_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i86_2_lut (.A(dec_new_block[85]), .B(round_key[85]), 
         .Z(block_new_127__N_1901[85])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i86_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i117_2_lut (.A(\block_reg[0] [20]), .B(round_key[116]), 
         .Z(\block_new_127__N_1645[116] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i117_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i85_2_lut (.A(dec_new_block[84]), .B(round_key[84]), 
         .Z(block_new_127__N_1901[84])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i85_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i116_2_lut (.A(\block_reg[0] [19]), .B(round_key[115]), 
         .Z(\block_new_127__N_1645[115] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i116_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i84_2_lut (.A(dec_new_block[83]), .B(round_key[83]), 
         .Z(block_new_127__N_1901[83])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i84_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i115_2_lut (.A(\block_reg[0] [18]), .B(round_key[114]), 
         .Z(\block_new_127__N_1645[114] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i115_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i83_2_lut (.A(dec_new_block[82]), .B(round_key[82]), 
         .Z(block_new_127__N_1901[82])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i83_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i114_2_lut (.A(\block_reg[0] [17]), .B(round_key[113]), 
         .Z(\block_new_127__N_1645[113] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i114_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i82_2_lut (.A(dec_new_block[81]), .B(round_key[81]), 
         .Z(block_new_127__N_1901[81])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i82_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i113_2_lut (.A(\block_reg[0] [16]), .B(round_key[112]), 
         .Z(block_new_127__N_1645_c[112])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i113_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i81_2_lut (.A(dec_new_block[80]), .B(round_key[80]), 
         .Z(block_new_127__N_1901[80])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i81_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i16_2_lut (.A(\block_reg[3] [15]), .B(round_key[15]), 
         .Z(block_new_127__N_1645_c[15])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i16_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i80_2_lut (.A(dec_new_block[79]), .B(round_key[79]), 
         .Z(block_new_127__N_1901[79])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i80_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i15_2_lut (.A(\block_reg[3] [14]), .B(round_key[14]), 
         .Z(\block_new_127__N_1645[14] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i15_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i79_2_lut (.A(dec_new_block[78]), .B(round_key[78]), 
         .Z(block_new_127__N_1901[78])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i79_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i14_2_lut (.A(\block_reg[3] [13]), .B(round_key[13]), 
         .Z(block_new_127__N_1645_c[13])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i14_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i78_2_lut (.A(dec_new_block[77]), .B(round_key[77]), 
         .Z(block_new_127__N_1901[77])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i78_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i13_2_lut (.A(\block_reg[3] [12]), .B(round_key[12]), 
         .Z(\block_new_127__N_1645[12] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i13_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i77_2_lut (.A(dec_new_block[76]), .B(round_key[76]), 
         .Z(block_new_127__N_1901[76])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i77_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i12_2_lut (.A(\block_reg[3] [11]), .B(round_key[11]), 
         .Z(block_new_127__N_1645_c[11])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i12_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i76_2_lut (.A(dec_new_block[75]), .B(round_key[75]), 
         .Z(block_new_127__N_1901[75])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i76_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i11_2_lut (.A(\block_reg[3] [10]), .B(round_key[10]), 
         .Z(\block_new_127__N_1645[10] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i11_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i75_2_lut (.A(dec_new_block[74]), .B(round_key[74]), 
         .Z(block_new_127__N_1901[74])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i75_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i10_2_lut (.A(\block_reg[3] [9]), .B(round_key[9]), 
         .Z(block_new_127__N_1645_c[9])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i10_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i74_2_lut (.A(dec_new_block[73]), .B(round_key[73]), 
         .Z(block_new_127__N_1901[73])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i74_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i9_2_lut (.A(\block_reg[3] [8]), .B(round_key[8]), 
         .Z(block_new_127__N_1645_c[8])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i9_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i73_2_lut (.A(dec_new_block[72]), .B(round_key[72]), 
         .Z(block_new_127__N_1901[72])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i73_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i40_2_lut (.A(\block_reg[2] [7]), .B(round_key[39]), 
         .Z(block_new_127__N_1645[39])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i40_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i72_2_lut (.A(dec_new_block[71]), .B(round_key[71]), 
         .Z(block_new_127__N_1901[71])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i72_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i39_2_lut (.A(\block_reg[2] [6]), .B(round_key[38]), 
         .Z(block_new_127__N_1645_c[38])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i39_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i71_2_lut (.A(dec_new_block[70]), .B(round_key[70]), 
         .Z(block_new_127__N_1901[70])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i71_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i38_2_lut (.A(\block_reg[2] [5]), .B(round_key[37]), 
         .Z(\block_new_127__N_1645[37] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i38_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i70_2_lut (.A(dec_new_block[69]), .B(round_key[69]), 
         .Z(block_new_127__N_1901[69])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i70_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i37_2_lut (.A(\block_reg[2] [4]), .B(round_key[36]), 
         .Z(\block_new_127__N_1645[36] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i37_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i69_2_lut (.A(dec_new_block[68]), .B(round_key[68]), 
         .Z(block_new_127__N_1901[68])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i69_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i36_2_lut (.A(\block_reg[2] [3]), .B(round_key[35]), 
         .Z(block_new_127__N_1645_c[35])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i36_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i68_2_lut (.A(dec_new_block[67]), .B(round_key[67]), 
         .Z(block_new_127__N_1901[67])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i68_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i35_2_lut (.A(\block_reg[2] [2]), .B(round_key[34]), 
         .Z(\block_new_127__N_1645[34] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i35_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i67_2_lut (.A(dec_new_block[66]), .B(round_key[66]), 
         .Z(block_new_127__N_1901[66])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i67_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i34_2_lut (.A(\block_reg[2] [1]), .B(round_key[33]), 
         .Z(\block_new_127__N_1645[33] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i34_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i66_2_lut (.A(dec_new_block[65]), .B(round_key[65]), 
         .Z(block_new_127__N_1901[65])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i66_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i33_2_lut (.A(\block_reg[2] [0]), .B(round_key[32]), 
         .Z(block_new_127__N_1645_c[32])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i33_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i65_2_lut (.A(dec_new_block[64]), .B(round_key[64]), 
         .Z(block_new_127__N_1901[64])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i65_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i64_2_lut (.A(\block_reg[2] [31]), .B(round_key[63]), 
         .Z(block_new_127__N_1645_c[63])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i64_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i64_2_lut (.A(dec_new_block[63]), .B(round_key[63]), 
         .Z(block_new_127__N_1901[63])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i64_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i63_2_lut (.A(\block_reg[2] [30]), .B(round_key[62]), 
         .Z(\block_new_127__N_1645[62] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i63_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i63_2_lut (.A(dec_new_block[62]), .B(round_key[62]), 
         .Z(block_new_127__N_1901[62])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i63_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i62_2_lut (.A(\block_reg[2] [29]), .B(round_key[61]), 
         .Z(\block_new_127__N_1645[61] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i62_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i62_2_lut (.A(dec_new_block[61]), .B(round_key[61]), 
         .Z(block_new_127__N_1901[61])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i62_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i61_2_lut (.A(\block_reg[2] [28]), .B(round_key[60]), 
         .Z(\block_new_127__N_1645[60] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i61_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i61_2_lut (.A(dec_new_block[60]), .B(round_key[60]), 
         .Z(block_new_127__N_1901[60])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i61_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i60_2_lut (.A(\block_reg[2] [27]), .B(round_key[59]), 
         .Z(\block_new_127__N_1645[59] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i60_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i60_2_lut (.A(dec_new_block[59]), .B(round_key[59]), 
         .Z(block_new_127__N_1901[59])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i60_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i59_2_lut (.A(\block_reg[2] [26]), .B(round_key[58]), 
         .Z(block_new_127__N_1645_c[58])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i59_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i59_2_lut (.A(dec_new_block[58]), .B(round_key[58]), 
         .Z(block_new_127__N_1901[58])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i59_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i58_2_lut (.A(\block_reg[2] [25]), .B(round_key[57]), 
         .Z(\block_new_127__N_1645[57] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i58_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i58_2_lut (.A(dec_new_block[57]), .B(round_key[57]), 
         .Z(block_new_127__N_1901[57])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i58_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i57_2_lut (.A(\block_reg[2] [24]), .B(round_key[56]), 
         .Z(block_new_127__N_1645_c[56])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i57_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i57_2_lut (.A(dec_new_block[56]), .B(round_key[56]), 
         .Z(block_new_127__N_1901[56])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i57_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i88_2_lut (.A(\block_reg[1] [23]), .B(round_key[87]), 
         .Z(\block_new_127__N_1645[87] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i88_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i56_2_lut (.A(dec_new_block[55]), .B(round_key[55]), 
         .Z(block_new_127__N_1901[55])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i56_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i87_2_lut (.A(\block_reg[1] [22]), .B(round_key[86]), 
         .Z(\block_new_127__N_1645[86] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i87_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i55_2_lut (.A(dec_new_block[54]), .B(round_key[54]), 
         .Z(block_new_127__N_1901[54])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i55_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i86_2_lut (.A(\block_reg[1] [21]), .B(round_key[85]), 
         .Z(\block_new_127__N_1645[85] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i86_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i54_2_lut (.A(dec_new_block[53]), .B(round_key[53]), 
         .Z(block_new_127__N_1901[53])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i54_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i85_2_lut (.A(\block_reg[1] [20]), .B(round_key[84]), 
         .Z(\block_new_127__N_1645[84] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i85_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i53_2_lut (.A(dec_new_block[52]), .B(round_key[52]), 
         .Z(block_new_127__N_1901[52])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i53_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i84_2_lut (.A(\block_reg[1] [19]), .B(round_key[83]), 
         .Z(\block_new_127__N_1645[83] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i84_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i52_2_lut (.A(dec_new_block[51]), .B(round_key[51]), 
         .Z(block_new_127__N_1901[51])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i52_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i83_2_lut (.A(\block_reg[1] [18]), .B(round_key[82]), 
         .Z(\block_new_127__N_1645[82] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i83_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i51_2_lut (.A(dec_new_block[50]), .B(round_key[50]), 
         .Z(block_new_127__N_1901[50])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i51_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i82_2_lut (.A(\block_reg[1] [17]), .B(round_key[81]), 
         .Z(\block_new_127__N_1645[81] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i82_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i50_2_lut (.A(dec_new_block[49]), .B(round_key[49]), 
         .Z(block_new_127__N_1901[49])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i50_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i81_2_lut (.A(\block_reg[1] [16]), .B(round_key[80]), 
         .Z(block_new_127__N_1645_c[80])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i81_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i49_2_lut (.A(dec_new_block[48]), .B(round_key[48]), 
         .Z(block_new_127__N_1901[48])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i49_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i112_2_lut (.A(\block_reg[0] [15]), .B(round_key[111]), 
         .Z(block_new_127__N_1645_c[111])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i112_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i48_2_lut (.A(dec_new_block[47]), .B(round_key[47]), 
         .Z(block_new_127__N_1901[47])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i48_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i111_2_lut (.A(\block_reg[0] [14]), .B(round_key[110]), 
         .Z(block_new_127__N_1645_c[110])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i111_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i47_2_lut (.A(dec_new_block[46]), .B(round_key[46]), 
         .Z(block_new_127__N_1901[46])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i47_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i110_2_lut (.A(\block_reg[0] [13]), .B(round_key[109]), 
         .Z(block_new_127__N_1645_c[109])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i110_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i46_2_lut (.A(dec_new_block[45]), .B(round_key[45]), 
         .Z(block_new_127__N_1901[45])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i46_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i109_2_lut (.A(\block_reg[0] [12]), .B(round_key[108]), 
         .Z(\block_new_127__N_1645[108] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i109_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i45_2_lut (.A(dec_new_block[44]), .B(round_key[44]), 
         .Z(block_new_127__N_1901[44])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i45_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i108_2_lut (.A(\block_reg[0] [11]), .B(round_key[107]), 
         .Z(\block_new_127__N_1645[107] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i108_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i44_2_lut (.A(dec_new_block[43]), .B(round_key[43]), 
         .Z(block_new_127__N_1901[43])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i44_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i107_2_lut (.A(\block_reg[0] [10]), .B(round_key[106]), 
         .Z(block_new_127__N_1645_c[106])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i107_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i43_2_lut (.A(dec_new_block[42]), .B(round_key[42]), 
         .Z(block_new_127__N_1901[42])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i43_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i106_2_lut (.A(\block_reg[0] [9]), .B(round_key[105]), 
         .Z(\block_new_127__N_1645[105] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i106_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i42_2_lut (.A(dec_new_block[41]), .B(round_key[41]), 
         .Z(block_new_127__N_1901[41])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i42_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i105_2_lut (.A(\block_reg[0] [8]), .B(round_key[104]), 
         .Z(block_new_127__N_1645_c[104])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i105_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i41_2_lut (.A(dec_new_block[40]), .B(round_key[40]), 
         .Z(block_new_127__N_1901[40])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i41_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i8_2_lut (.A(\block_reg[3] [7]), .B(round_key[7]), 
         .Z(\block_new_127__N_1645[7] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i8_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i40_2_lut (.A(dec_new_block[39]), .B(round_key[39]), 
         .Z(block_new_127__N_1901[39])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i40_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i7_2_lut (.A(\block_reg[3] [6]), .B(round_key[6]), 
         .Z(block_new_127__N_1645_c[6])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i7_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i39_2_lut (.A(dec_new_block[38]), .B(round_key[38]), 
         .Z(block_new_127__N_1901[38])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i39_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i6_2_lut (.A(\block_reg[3] [5]), .B(round_key[5]), 
         .Z(\block_new_127__N_1645[5] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i6_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i38_2_lut (.A(dec_new_block[37]), .B(round_key[37]), 
         .Z(block_new_127__N_1901[37])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i38_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i5_2_lut (.A(\block_reg[3] [4]), .B(round_key[4]), 
         .Z(\block_new_127__N_1645[4] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i5_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i37_2_lut (.A(dec_new_block[36]), .B(round_key[36]), 
         .Z(block_new_127__N_1901[36])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i37_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i4_2_lut (.A(\block_reg[3] [3]), .B(round_key[3]), 
         .Z(\block_new_127__N_1645[3] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i4_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i36_2_lut (.A(dec_new_block[35]), .B(round_key[35]), 
         .Z(block_new_127__N_1901[35])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i36_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i3_2_lut (.A(\block_reg[3] [2]), .B(round_key[2]), 
         .Z(\block_new_127__N_1645[2] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i3_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i35_2_lut (.A(dec_new_block[34]), .B(round_key[34]), 
         .Z(block_new_127__N_1901[34])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i35_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i2_2_lut (.A(\block_reg[3] [1]), .B(round_key[1]), 
         .Z(\block_new_127__N_1645[1] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i2_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i34_2_lut (.A(dec_new_block[33]), .B(round_key[33]), 
         .Z(block_new_127__N_1901[33])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i34_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i1_2_lut (.A(\block_reg[3] [0]), .B(round_key[0]), 
         .Z(block_new_127__N_1645_c[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i1_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i33_2_lut (.A(dec_new_block[32]), .B(round_key[32]), 
         .Z(block_new_127__N_1901[32])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i33_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i32_2_lut (.A(\block_reg[3] [31]), .B(round_key[31]), 
         .Z(block_new_127__N_1645_c[31])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i32_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i32_2_lut (.A(dec_new_block[31]), .B(round_key[31]), 
         .Z(block_new_127__N_1901[31])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i32_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i31_2_lut (.A(\block_reg[3] [30]), .B(round_key[30]), 
         .Z(\block_new_127__N_1645[30] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i31_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i31_2_lut (.A(dec_new_block[30]), .B(round_key[30]), 
         .Z(block_new_127__N_1901[30])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i31_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i30_2_lut (.A(\block_reg[3] [29]), .B(round_key[29]), 
         .Z(block_new_127__N_1645_c[29])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i30_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i30_2_lut (.A(dec_new_block[29]), .B(round_key[29]), 
         .Z(block_new_127__N_1901[29])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i30_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i29_2_lut (.A(\block_reg[3] [28]), .B(round_key[28]), 
         .Z(\block_new_127__N_1645[28] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i29_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i29_2_lut (.A(dec_new_block[28]), .B(round_key[28]), 
         .Z(block_new_127__N_1901[28])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i29_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i28_2_lut (.A(\block_reg[3] [27]), .B(round_key[27]), 
         .Z(\block_new_127__N_1645[27] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i28_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i28_2_lut (.A(dec_new_block[27]), .B(round_key[27]), 
         .Z(block_new_127__N_1901[27])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i28_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i27_2_lut (.A(\block_reg[3] [26]), .B(round_key[26]), 
         .Z(block_new_127__N_1645_c[26])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i27_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i27_2_lut (.A(dec_new_block[26]), .B(round_key[26]), 
         .Z(block_new_127__N_1901[26])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i27_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i26_2_lut (.A(\block_reg[3] [25]), .B(round_key[25]), 
         .Z(\block_new_127__N_1645[25] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i26_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i26_2_lut (.A(dec_new_block[25]), .B(round_key[25]), 
         .Z(block_new_127__N_1901[25])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i26_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i25_2_lut (.A(\block_reg[3] [24]), .B(round_key[24]), 
         .Z(block_new_127__N_1645_c[24])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i25_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i25_2_lut (.A(dec_new_block[24]), .B(round_key[24]), 
         .Z(block_new_127__N_1901[24])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i25_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i56_2_lut (.A(\block_reg[2] [23]), .B(round_key[55]), 
         .Z(block_new_127__N_1645_c[55])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i56_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i24_2_lut (.A(dec_new_block[23]), .B(round_key[23]), 
         .Z(block_new_127__N_1901[23])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i24_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i55_2_lut (.A(\block_reg[2] [22]), .B(round_key[54]), 
         .Z(block_new_127__N_1645_c[54])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i55_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i23_2_lut (.A(dec_new_block[22]), .B(round_key[22]), 
         .Z(block_new_127__N_1901[22])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i23_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i54_2_lut (.A(\block_reg[2] [21]), .B(round_key[53]), 
         .Z(block_new_127__N_1645_c[53])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i54_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i22_2_lut (.A(dec_new_block[21]), .B(round_key[21]), 
         .Z(block_new_127__N_1901[21])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i22_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i53_2_lut (.A(\block_reg[2] [20]), .B(round_key[52]), 
         .Z(block_new_127__N_1645_c[52])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i53_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i21_2_lut (.A(dec_new_block[20]), .B(round_key[20]), 
         .Z(block_new_127__N_1901[20])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i21_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i52_2_lut (.A(\block_reg[2] [19]), .B(round_key[51]), 
         .Z(\block_new_127__N_1645[51] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i52_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i20_2_lut (.A(dec_new_block[19]), .B(round_key[19]), 
         .Z(block_new_127__N_1901[19])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i20_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i51_2_lut (.A(\block_reg[2] [18]), .B(round_key[50]), 
         .Z(\block_new_127__N_1645[50] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i51_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i19_2_lut (.A(dec_new_block[18]), .B(round_key[18]), 
         .Z(block_new_127__N_1901[18])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i19_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i50_2_lut (.A(\block_reg[2] [17]), .B(round_key[49]), 
         .Z(\block_new_127__N_1645[49] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i50_2_lut.init = 16'h6666;
    LUT4 i3_2_lut_3_lut_4_lut_adj_230 (.A(block_new_127__N_1901[57]), .B(block_new_127__N_1901[49]), 
         .C(n33810), .D(n33811), .Z(n9_adj_8010)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i3_2_lut_3_lut_4_lut_adj_230.init = 16'h6996;
    LUT4 new_block_127__I_0_i18_2_lut (.A(dec_new_block[17]), .B(round_key[17]), 
         .Z(block_new_127__N_1901[17])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i18_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i49_2_lut (.A(\block_reg[2] [16]), .B(round_key[48]), 
         .Z(block_new_127__N_1645_c[48])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i49_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i17_2_lut (.A(dec_new_block[16]), .B(round_key[16]), 
         .Z(block_new_127__N_1901[16])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i17_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i80_2_lut (.A(\block_reg[1] [15]), .B(round_key[79]), 
         .Z(block_new_127__N_1645_c[79])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i80_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i16_2_lut (.A(dec_new_block[15]), .B(round_key[15]), 
         .Z(block_new_127__N_1901[15])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i16_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i79_2_lut (.A(\block_reg[1] [14]), .B(round_key[78]), 
         .Z(block_new_127__N_1645_c[78])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i79_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i15_2_lut (.A(dec_new_block[14]), .B(round_key[14]), 
         .Z(block_new_127__N_1901[14])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i15_2_lut.init = 16'h6666;
    LUT4 i2_3_lut_4_lut_adj_231 (.A(n33788), .B(n33778), .C(n12810), .D(n33697), 
         .Z(n29273)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i2_3_lut_4_lut_adj_231.init = 16'h6996;
    LUT4 i1_2_lut_3_lut_adj_232 (.A(block_new_127__N_1901[63]), .B(block_new_127__N_1901[56]), 
         .C(block_new_127__N_1901[48]), .Z(n4_adj_7932)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_3_lut_adj_232.init = 16'h9696;
    LUT4 block_127__I_0_i78_2_lut (.A(\block_reg[1] [13]), .B(round_key[77]), 
         .Z(block_new_127__N_1645_c[77])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i78_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i14_2_lut (.A(dec_new_block[13]), .B(round_key[13]), 
         .Z(block_new_127__N_1901[13])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i14_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i77_2_lut (.A(\block_reg[1] [12]), .B(round_key[76]), 
         .Z(\block_new_127__N_1645[76] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i77_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i13_2_lut (.A(dec_new_block[12]), .B(round_key[12]), 
         .Z(block_new_127__N_1901[12])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i13_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i76_2_lut (.A(\block_reg[1] [11]), .B(round_key[75]), 
         .Z(\block_new_127__N_1645[75] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i76_2_lut.init = 16'h6666;
    LUT4 i1_2_lut_rep_408_3_lut_4_lut (.A(block_new_127__N_1901[37]), .B(block_new_127__N_1901[32]), 
         .C(block_new_127__N_1901[56]), .D(block_new_127__N_1901[63]), .Z(n33712)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_408_3_lut_4_lut.init = 16'h6996;
    LUT4 new_block_127__I_0_i12_2_lut (.A(dec_new_block[11]), .B(round_key[11]), 
         .Z(block_new_127__N_1901[11])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i12_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i75_2_lut (.A(\block_reg[1] [10]), .B(round_key[74]), 
         .Z(block_new_127__N_1645_c[74])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i75_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i11_2_lut (.A(dec_new_block[10]), .B(round_key[10]), 
         .Z(block_new_127__N_1901[10])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i11_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i74_2_lut (.A(\block_reg[1] [9]), .B(round_key[73]), 
         .Z(\block_new_127__N_1645[73] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i74_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i10_2_lut (.A(dec_new_block[9]), .B(round_key[9]), 
         .Z(block_new_127__N_1901[9])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i10_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i73_2_lut (.A(\block_reg[1] [8]), .B(round_key[72]), 
         .Z(block_new_127__N_1645_c[72])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i73_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i9_2_lut (.A(dec_new_block[8]), .B(round_key[8]), 
         .Z(block_new_127__N_1901[8])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i9_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i104_2_lut (.A(\block_reg[0] [7]), .B(round_key[103]), 
         .Z(block_new_127__N_1645_c[103])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i104_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i8_2_lut (.A(dec_new_block[7]), .B(round_key[7]), 
         .Z(block_new_127__N_1901[7])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i8_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i103_2_lut (.A(\block_reg[0] [6]), .B(round_key[102]), 
         .Z(\block_new_127__N_1645[102] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i103_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i7_2_lut (.A(dec_new_block[6]), .B(round_key[6]), 
         .Z(block_new_127__N_1901[6])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i7_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i102_2_lut (.A(\block_reg[0] [5]), .B(round_key[101]), 
         .Z(block_new_127__N_1645_c[101])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i102_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i126_2_lut (.A(\block_reg[0] [29]), .B(round_key[125]), 
         .Z(\block_new_127__N_1645[125] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i126_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i6_2_lut (.A(dec_new_block[5]), .B(round_key[5]), 
         .Z(block_new_127__N_1901[5])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i6_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i101_2_lut (.A(\block_reg[0] [4]), .B(round_key[100]), 
         .Z(block_new_127__N_1645_c[100])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i101_2_lut.init = 16'h6666;
    LUT4 i1_4_lut_adj_233 (.A(n14912), .B(n149), .C(n14919), .D(n110), 
         .Z(n152)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(96[7:17])
    defparam i1_4_lut_adj_233.init = 16'hc088;
    LUT4 new_block_127__I_0_i5_2_lut (.A(dec_new_block[4]), .B(round_key[4]), 
         .Z(block_new_127__N_1901[4])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i5_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i100_2_lut (.A(\block_reg[0] [3]), .B(round_key[99]), 
         .Z(\block_new_127__N_1645[99] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i100_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i4_2_lut (.A(dec_new_block[3]), .B(round_key[3]), 
         .Z(block_new_127__N_1901[3])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i4_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i99_2_lut (.A(\block_reg[0] [2]), .B(round_key[98]), 
         .Z(\block_new_127__N_1645[98] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i99_2_lut.init = 16'h6666;
    LUT4 new_block_127__I_0_i3_2_lut (.A(dec_new_block[2]), .B(round_key[2]), 
         .Z(block_new_127__N_1901[2])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i3_2_lut.init = 16'h6666;
    LUT4 block_127__I_0_i98_2_lut (.A(\block_reg[0] [1]), .B(round_key[97]), 
         .Z(\block_new_127__N_1645[97] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i98_2_lut.init = 16'h6666;
    LUT4 i4_3_lut_4_lut_adj_234 (.A(n33788), .B(n33778), .C(block_new_127__N_1901[22]), 
         .D(block_new_127__N_1901[29]), .Z(n10_adj_7818)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i4_3_lut_4_lut_adj_234.init = 16'h6996;
    LUT4 new_block_127__I_0_i126_2_lut (.A(dec_new_block[125]), .B(round_key[125]), 
         .Z(block_new_127__N_1901[125])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i126_2_lut.init = 16'h6666;
    LUT4 i3_2_lut_3_lut_4_lut_adj_235 (.A(block_new_127__N_1901[37]), .B(block_new_127__N_1901[32]), 
         .C(n29471), .D(block_new_127__N_1901[40]), .Z(n9_adj_7833)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i3_2_lut_3_lut_4_lut_adj_235.init = 16'h6996;
    LUT4 i2_2_lut_3_lut_4_lut_adj_236 (.A(block_new_127__N_1901[37]), .B(block_new_127__N_1901[32]), 
         .C(block_new_127__N_1901[63]), .D(block_new_127__N_1901[40]), .Z(n7_adj_7727)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i2_2_lut_3_lut_4_lut_adj_236.init = 16'h6996;
    LUT4 i1_2_lut_3_lut_4_lut_adj_237 (.A(block_new_127__N_1901[37]), .B(block_new_127__N_1901[32]), 
         .C(n33812), .D(block_new_127__N_1901[39]), .Z(n5_adj_7771)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_3_lut_4_lut_adj_237.init = 16'h6996;
    LUT4 i3_3_lut_4_lut_adj_238 (.A(block_new_127__N_1901[47]), .B(block_new_127__N_1901[55]), 
         .C(n12071), .D(n33812), .Z(n29471)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i3_3_lut_4_lut_adj_238.init = 16'h6996;
    LUT4 i1_2_lut_3_lut_adj_239 (.A(block_new_127__N_1901[47]), .B(block_new_127__N_1901[55]), 
         .C(block_new_127__N_1901[63]), .Z(n5_adj_7742)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_3_lut_adj_239.init = 16'h9696;
    LUT4 new_block_127__I_0_i2_2_lut (.A(dec_new_block[1]), .B(round_key[1]), 
         .Z(block_new_127__N_1901[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i2_2_lut.init = 16'h6666;
    LUT4 i1_2_lut_3_lut_4_lut_adj_240 (.A(block_new_127__N_1901[47]), .B(block_new_127__N_1901[55]), 
         .C(block_new_127__N_1901[54]), .D(block_new_127__N_1901[62]), .Z(n4_adj_7738)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_3_lut_4_lut_adj_240.init = 16'h6996;
    LUT4 i176_3_lut (.A(n6363[0]), .B(n6363[2]), .C(n33856), .Z(n2886)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(221[17:29])
    defparam i176_3_lut.init = 16'hecec;
    LUT4 i1_2_lut_rep_381_3_lut (.A(block_new_127__N_1901[45]), .B(block_new_127__N_1901[61]), 
         .C(block_new_127__N_1901[39]), .Z(n33685)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_rep_381_3_lut.init = 16'h9696;
    LUT4 i2_2_lut_3_lut_4_lut_adj_241 (.A(block_new_127__N_1901[45]), .B(block_new_127__N_1901[61]), 
         .C(block_new_127__N_1901[40]), .D(block_new_127__N_1901[37]), .Z(n6_adj_8018)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i2_2_lut_3_lut_4_lut_adj_241.init = 16'h6996;
    LUT4 i1_2_lut_rep_407_3_lut (.A(block_new_127__N_1901[45]), .B(block_new_127__N_1901[61]), 
         .C(block_new_127__N_1901[37]), .Z(n33711)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_rep_407_3_lut.init = 16'h9696;
    LUT4 i1_4_lut_adj_242 (.A(n14890), .B(n6362[3]), .C(n166), .D(n6363[1]), 
         .Z(n28836)) /* synthesis lut_function=(A+(B (C)+!B (C+(D)))) */ ;
    defparam i1_4_lut_adj_242.init = 16'hfbfa;
    LUT4 i178_3_lut (.A(encdec_reg), .B(dec_ctrl_new_2__N_2032), .C(\aes_core_ctrl_new_1__N_858[1] ), 
         .Z(n166)) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes.v(96[7:17])
    defparam i178_3_lut.init = 16'h8c8c;
    LUT4 mux_626_Mux_7_i2_4_lut (.A(new_sboxw[7]), .B(n11_adj_8017), .C(update_type[0]), 
         .D(n12_adj_8003), .Z(n2_adj_8019)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(319[7] 388[14])
    defparam mux_626_Mux_7_i2_4_lut.init = 16'h3aca;
    LUT4 i3_3_lut_4_lut_adj_243 (.A(n33788), .B(n33778), .C(block_new_127__N_1901[6]), 
         .D(n33827), .Z(n8_adj_7875)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i3_3_lut_4_lut_adj_243.init = 16'h6996;
    LUT4 i2_2_lut_3_lut_4_lut_adj_244 (.A(block_new_127__N_1901[39]), .B(block_new_127__N_1901[40]), 
         .C(n29393), .D(block_new_127__N_1901[57]), .Z(n6_adj_8008)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i2_2_lut_3_lut_4_lut_adj_244.init = 16'h6996;
    LUT4 i2_2_lut_3_lut_adj_245 (.A(block_new_127__N_1901[42]), .B(block_new_127__N_1901[47]), 
         .C(block_new_127__N_1901[59]), .Z(n7_adj_7975)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i2_2_lut_3_lut_adj_245.init = 16'h9696;
    LUT4 block_127__I_0_i97_2_lut (.A(\block_reg[0] [0]), .B(round_key[96]), 
         .Z(block_new_127__N_1645_c[96])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam block_127__I_0_i97_2_lut.init = 16'h6666;
    LUT4 i1_2_lut_3_lut_adj_246 (.A(block_new_127__N_1901[42]), .B(block_new_127__N_1901[47]), 
         .C(n11890), .Z(n5_adj_7901)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_3_lut_adj_246.init = 16'h9696;
    LUT4 i2_2_lut_3_lut_4_lut_adj_247 (.A(block_new_127__N_1901[126]), .B(n33766), 
         .C(n33759), .D(block_new_127__N_1901[106]), .Z(n7_adj_7753)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i2_2_lut_3_lut_4_lut_adj_247.init = 16'h6996;
    LUT4 i1_4_lut_adj_248 (.A(block_new_127__N_1901[109]), .B(n33715), .C(n33714), 
         .D(block_new_127__N_1901[118]), .Z(n29160)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_4_lut_adj_248.init = 16'h6996;
    LUT4 i1_4_lut_adj_249 (.A(dec_ctrl_new_2__N_2032), .B(n33842), .C(n20702), 
         .D(n33844), .Z(block_w2_we)) /* synthesis lut_function=(!(A+!(B (C+(D))+!B !((D)+!C)))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(462[7] 518[14])
    defparam i1_4_lut_adj_249.init = 16'h4450;
    LUT4 i4_4_lut_adj_250 (.A(n12084), .B(n29429), .C(n29375), .D(n6_adj_8020), 
         .Z(n28961)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i4_4_lut_adj_250.init = 16'h6996;
    LUT4 i1_4_lut_adj_251 (.A(block_new_127__N_1901[113]), .B(block_new_127__N_1901[97]), 
         .C(block_new_127__N_1901[118]), .D(block_new_127__N_1901[102]), 
         .Z(n29220)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_4_lut_adj_251.init = 16'h6996;
    LUT4 i3_3_lut_4_lut_adj_252 (.A(block_new_127__N_1901[113]), .B(n33767), 
         .C(n33768), .D(n33518), .Z(n8_adj_7878)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i3_3_lut_4_lut_adj_252.init = 16'h6996;
    LUT4 xor_638_i5_2_lut_3_lut (.A(block_new_127__N_1901[17]), .B(block_new_127__N_1901[22]), 
         .C(block_new_127__N_1901[21]), .Z(n6111[4])) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam xor_638_i5_2_lut_3_lut.init = 16'h9696;
    LUT4 i5_4_lut_adj_253 (.A(n9_adj_8021), .B(block_new_127__N_1901[29]), 
         .C(n8_adj_8022), .D(n6345[3]), .Z(n29447)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i5_4_lut_adj_253.init = 16'h6996;
    LUT4 i2_2_lut_3_lut_4_lut_adj_254 (.A(n33837), .B(n33838), .C(n33710), 
         .D(block_new_127__N_1901[101]), .Z(n6_adj_7720)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i2_2_lut_3_lut_4_lut_adj_254.init = 16'h6996;
    LUT4 i2_3_lut (.A(block_new_127__N_1901[0]), .B(block_new_127__N_1901[7]), 
         .C(block_new_127__N_1901[5]), .Z(n6345[3])) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i2_3_lut.init = 16'h9696;
    LUT4 i1_2_lut_3_lut_adj_255 (.A(block_new_127__N_1901[66]), .B(block_new_127__N_1901[71]), 
         .C(block_new_127__N_1901[91]), .Z(n29172)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_3_lut_adj_255.init = 16'h9696;
    LUT4 i1_2_lut_3_lut_4_lut_adj_256 (.A(block_new_127__N_1901[124]), .B(n33770), 
         .C(n33766), .D(block_new_127__N_1901[126]), .Z(n5_adj_7719)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_3_lut_4_lut_adj_256.init = 16'h6996;
    LUT4 i1_2_lut_3_lut_4_lut_adj_257 (.A(block_new_127__N_1901[92]), .B(n33797), 
         .C(n33704), .D(block_new_127__N_1901[84]), .Z(n5_adj_7896)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_3_lut_4_lut_adj_257.init = 16'h6996;
    LUT4 i4_4_lut_adj_258 (.A(n33522), .B(block_new_127__N_1901[91]), .C(block_new_127__N_1901[75]), 
         .D(n33822), .Z(n10_adj_7988)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i4_4_lut_adj_258.init = 16'h6996;
    LUT4 i2_2_lut_3_lut_adj_259 (.A(block_new_127__N_1901[18]), .B(block_new_127__N_1901[23]), 
         .C(block_new_127__N_1901[19]), .Z(n7_adj_7984)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i2_2_lut_3_lut_adj_259.init = 16'h9696;
    LUT4 i2_2_lut_3_lut_adj_260 (.A(block_new_127__N_1901[18]), .B(block_new_127__N_1901[23]), 
         .C(n29181), .Z(n6_adj_7979)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i2_2_lut_3_lut_adj_260.init = 16'h9696;
    LUT4 i2_2_lut_4_lut_adj_261 (.A(n29480), .B(block_new_127__N_1901[59]), 
         .C(block_new_127__N_1901[43]), .D(n33806), .Z(n6_adj_7902)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i2_2_lut_4_lut_adj_261.init = 16'h6996;
    LUT4 i1_2_lut_3_lut_adj_262 (.A(block_new_127__N_1901[26]), .B(block_new_127__N_1901[31]), 
         .C(n29181), .Z(n5_adj_7915)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_3_lut_adj_262.init = 16'h9696;
    LUT4 i1_4_lut_adj_263 (.A(block_new_127__N_1901[65]), .B(block_new_127__N_1901[81]), 
         .C(block_new_127__N_1901[70]), .D(block_new_127__N_1901[86]), .Z(n29199)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_4_lut_adj_263.init = 16'h6996;
    LUT4 i4_4_lut_adj_264 (.A(n12074), .B(n29432), .C(n33819), .D(n6_adj_8023), 
         .Z(n29254)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i4_4_lut_adj_264.init = 16'h6996;
    LUT4 i3_3_lut_4_lut_adj_265 (.A(block_new_127__N_1901[26]), .B(block_new_127__N_1901[31]), 
         .C(block_new_127__N_1901[11]), .D(n33508), .Z(n8_adj_7985)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i3_3_lut_4_lut_adj_265.init = 16'h6996;
    LUT4 i2_2_lut_3_lut_adj_266 (.A(block_new_127__N_1901[87]), .B(block_new_127__N_1901[80]), 
         .C(block_new_127__N_1901[64]), .Z(n7_adj_7850)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i2_2_lut_3_lut_adj_266.init = 16'h9696;
    LUT4 i2_3_lut_adj_267 (.A(block_new_127__N_1901[88]), .B(block_new_127__N_1901[95]), 
         .C(block_new_127__N_1901[93]), .Z(n3564[3])) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i2_3_lut_adj_267.init = 16'h9696;
    LUT4 i2_3_lut_adj_268 (.A(block_new_127__N_1901[85]), .B(block_new_127__N_1901[77]), 
         .C(block_new_127__N_1901[69]), .Z(n29432)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i2_3_lut_adj_268.init = 16'h9696;
    LUT4 i1_2_lut_3_lut_adj_269 (.A(block_new_127__N_1901[79]), .B(block_new_127__N_1901[72]), 
         .C(n3564[3]), .Z(n6_adj_8023)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_3_lut_adj_269.init = 16'h9696;
    LUT4 i1_4_lut_adj_270 (.A(block_new_127__N_1901[89]), .B(block_new_127__N_1901[73]), 
         .C(block_new_127__N_1901[94]), .D(block_new_127__N_1901[78]), .Z(n29483)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_4_lut_adj_270.init = 16'h6996;
    LUT4 i3_4_lut (.A(block_new_127__N_1901[27]), .B(block_new_127__N_1901[11]), 
         .C(n33815), .D(n6327[3]), .Z(n29181)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i3_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_4_lut_adj_271 (.A(n33784), .B(n33817), .C(n33823), .D(block_new_127__N_1901[28]), 
         .Z(n5_adj_7918)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_4_lut_adj_271.init = 16'h6996;
    LUT4 i3_4_lut_adj_272 (.A(block_new_127__N_1901[35]), .B(n33712), .C(n33813), 
         .D(n29471), .Z(n11890)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i3_4_lut_adj_272.init = 16'h6996;
    LUT4 i1_4_lut_adj_273 (.A(block_new_127__N_1901[41]), .B(block_new_127__N_1901[57]), 
         .C(block_new_127__N_1901[46]), .D(block_new_127__N_1901[62]), .Z(n29408)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_4_lut_adj_273.init = 16'h6996;
    LUT4 i1_2_lut_4_lut_adj_274 (.A(n33784), .B(n33817), .C(n33823), .D(n11918), 
         .Z(n4_adj_7869)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_4_lut_adj_274.init = 16'h6996;
    LUT4 i3_2_lut_3_lut_adj_275 (.A(block_new_127__N_1901[82]), .B(block_new_127__N_1901[87]), 
         .C(n29199), .Z(n9_adj_7987)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i3_2_lut_3_lut_adj_275.init = 16'h9696;
    LUT4 i2_3_lut_rep_281_4_lut (.A(block_new_127__N_1901[37]), .B(n33798), 
         .C(n4770[4]), .D(block_new_127__N_1901[45]), .Z(n33585)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i2_3_lut_rep_281_4_lut.init = 16'h6996;
    LUT4 i1_4_lut_adj_276 (.A(block_new_127__N_1901[38]), .B(block_new_127__N_1901[54]), 
         .C(n6_adj_8018), .D(block_new_127__N_1901[53]), .Z(n28926)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_4_lut_adj_276.init = 16'h6996;
    LUT4 i1_2_lut_3_lut_adj_277 (.A(block_new_127__N_1901[74]), .B(block_new_127__N_1901[79]), 
         .C(block_new_127__N_1901[83]), .Z(n5_adj_7982)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_3_lut_adj_277.init = 16'h9696;
    LUT4 i2_2_lut_3_lut_4_lut_adj_278 (.A(block_new_127__N_1901[2]), .B(block_new_127__N_1901[7]), 
         .C(n29447), .D(block_new_127__N_1901[19]), .Z(n6_adj_7916)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i2_2_lut_3_lut_4_lut_adj_278.init = 16'h6996;
    LUT4 i1_2_lut_rep_282_4_lut (.A(n5085[3]), .B(n33786), .C(n33806), 
         .D(n33706), .Z(n33586)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_rep_282_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_409_3_lut (.A(block_new_127__N_1901[2]), .B(block_new_127__N_1901[7]), 
         .C(block_new_127__N_1901[19]), .Z(n33713)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_rep_409_3_lut.init = 16'h9696;
    LUT4 i1_2_lut_4_lut_adj_279 (.A(n5085[3]), .B(n33786), .C(n33806), 
         .D(n12921), .Z(n5_adj_7799)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_4_lut_adj_279.init = 16'h6996;
    LUT4 i4_4_lut_adj_280 (.A(n7_adj_8005), .B(n29480), .C(block_new_127__N_1901[45]), 
         .D(block_new_127__N_1901[37]), .Z(n12921)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i4_4_lut_adj_280.init = 16'h6996;
    LUT4 i1_2_lut_3_lut_adj_281 (.A(block_new_127__N_1901[10]), .B(block_new_127__N_1901[15]), 
         .C(block_new_127__N_1901[27]), .Z(n5_adj_7990)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_3_lut_adj_281.init = 16'h9696;
    LUT4 i1_4_lut_adj_282 (.A(block_new_127__N_1901[49]), .B(block_new_127__N_1901[33]), 
         .C(block_new_127__N_1901[54]), .D(block_new_127__N_1901[38]), .Z(n29480)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_4_lut_adj_282.init = 16'h6996;
    LUT4 new_block_127__I_0_i128_2_lut (.A(dec_new_block[127]), .B(round_key[127]), 
         .Z(block_new_127__N_1901[127])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(186[21:32])
    defparam new_block_127__I_0_i128_2_lut.init = 16'h6666;
    LUT4 i1_2_lut_3_lut_4_lut_adj_283 (.A(block_new_127__N_1901[10]), .B(block_new_127__N_1901[15]), 
         .C(n29447), .D(block_new_127__N_1901[3]), .Z(n5_adj_7978)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_3_lut_4_lut_adj_283.init = 16'h6996;
    LUT4 i2_2_lut_3_lut_4_lut_adj_284 (.A(block_new_127__N_1901[15]), .B(block_new_127__N_1901[8]), 
         .C(block_new_127__N_1901[24]), .D(block_new_127__N_1901[31]), .Z(n8_adj_8022)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i2_2_lut_3_lut_4_lut_adj_284.init = 16'h6996;
    LUT4 i1_2_lut_3_lut_4_lut_adj_285 (.A(block_new_127__N_1901[60]), .B(n33787), 
         .C(n33799), .D(block_new_127__N_1901[44]), .Z(n5_adj_7774)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_3_lut_4_lut_adj_285.init = 16'h6996;
    LUT4 i3_4_lut_adj_286 (.A(block_new_127__N_1901[93]), .B(n29432), .C(n29199), 
         .D(n29483), .Z(n12748)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i3_4_lut_adj_286.init = 16'h6996;
    LUT4 i2_2_lut (.A(n29199), .B(n29254), .Z(n6_adj_7947)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i2_2_lut.init = 16'h6666;
    LUT4 i2_2_lut_3_lut_4_lut_adj_287 (.A(block_new_127__N_1901[60]), .B(n33787), 
         .C(n33763), .D(n33798), .Z(n6_adj_7800)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i2_2_lut_3_lut_4_lut_adj_287.init = 16'h6996;
    LUT4 i3_2_lut_3_lut_4_lut_adj_288 (.A(block_new_127__N_1901[23]), .B(block_new_127__N_1901[16]), 
         .C(block_new_127__N_1901[13]), .D(block_new_127__N_1901[21]), .Z(n9_adj_8021)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i3_2_lut_3_lut_4_lut_adj_288.init = 16'h6996;
    LUT4 i3_4_lut_adj_289 (.A(n33791), .B(n873[3]), .C(n648[3]), .D(n29220), 
         .Z(n29444)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i3_4_lut_adj_289.init = 16'h6996;
    LUT4 i2_2_lut_3_lut_4_lut_adj_290 (.A(block_new_127__N_1901[100]), .B(n33838), 
         .C(n33715), .D(n33790), .Z(n6_adj_7939)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i2_2_lut_3_lut_4_lut_adj_290.init = 16'h6996;
    LUT4 i3_4_lut_adj_291 (.A(n33788), .B(n6111[4]), .C(n8_adj_8000), 
         .D(n6048[4]), .Z(n29288)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i3_4_lut_adj_291.init = 16'h6996;
    LUT4 i3_4_lut_adj_292 (.A(n33818), .B(block_new_127__N_1901[30]), .C(n33824), 
         .D(block_new_127__N_1901[14]), .Z(n12810)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i3_4_lut_adj_292.init = 16'h6996;
    LUT4 xor_631_i5_2_lut_3_lut (.A(block_new_127__N_1901[25]), .B(block_new_127__N_1901[30]), 
         .C(block_new_127__N_1901[29]), .Z(n6048[4])) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam xor_631_i5_2_lut_3_lut.init = 16'h9696;
    LUT4 i1_2_lut_4_lut_adj_293 (.A(n33795), .B(n33822), .C(n33809), .D(block_new_127__N_1901[92]), 
         .Z(n5_adj_7952)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_4_lut_adj_293.init = 16'h6996;
    LUT4 i3_4_lut_adj_294 (.A(block_new_127__N_1901[4]), .B(n8_adj_8000), 
         .C(n6111[4]), .D(n6048[4]), .Z(n29291)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i3_4_lut_adj_294.init = 16'h6996;
    LUT4 i1_2_lut_rep_216_4_lut (.A(n33801), .B(n33805), .C(n33814), .D(n12921), 
         .Z(n33520)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i1_2_lut_rep_216_4_lut.init = 16'h6996;
    LUT4 i4_4_lut_adj_295 (.A(n33695), .B(n33775), .C(block_new_127__N_1901[2]), 
         .D(n6_adj_7999), .Z(n28882)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i4_4_lut_adj_295.init = 16'h6996;
    LUT4 i2_2_lut_3_lut_4_lut_adj_296 (.A(n33799), .B(n33798), .C(n12921), 
         .D(n33706), .Z(n6_adj_7956)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i2_2_lut_3_lut_4_lut_adj_296.init = 16'h6996;
    LUT4 i1_2_lut_4_lut_adj_297 (.A(block_new_127__N_1901[115]), .B(n33834), 
         .C(block_new_127__N_1901[123]), .D(n33833), .Z(n4_adj_7961)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_4_lut_adj_297.init = 16'h6996;
    LUT4 i3_4_lut_adj_298 (.A(n33839), .B(block_new_127__N_1901[119]), .C(n33691), 
         .D(block_new_127__N_1901[103]), .Z(n29231)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i3_4_lut_adj_298.init = 16'h6996;
    LUT4 i2_2_lut_4_lut_adj_299 (.A(block_new_127__N_1901[115]), .B(n33834), 
         .C(block_new_127__N_1901[123]), .D(n28961), .Z(n7_adj_7888)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i2_2_lut_4_lut_adj_299.init = 16'h6996;
    LUT4 i1_3_lut_4_lut (.A(block_new_127__N_1901[109]), .B(block_new_127__N_1901[111]), 
         .C(block_new_127__N_1901[104]), .D(block_new_127__N_1901[96]), 
         .Z(n29375)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_3_lut_4_lut.init = 16'h6996;
    LUT4 i2_2_lut_3_lut_4_lut_adj_300 (.A(block_new_127__N_1901[71]), .B(n33803), 
         .C(n33796), .D(block_new_127__N_1901[88]), .Z(n6_adj_7762)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i2_2_lut_3_lut_4_lut_adj_300.init = 16'h6996;
    LUT4 i3_4_lut_adj_301 (.A(block_new_127__N_1901[14]), .B(n33789), .C(block_new_127__N_1901[20]), 
         .D(n33687), .Z(n29143)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i3_4_lut_adj_301.init = 16'h6996;
    LUT4 i2_3_lut_rep_286_4_lut (.A(block_new_127__N_1901[71]), .B(n33803), 
         .C(block_new_127__N_1901[94]), .D(block_new_127__N_1901[79]), .Z(n33590)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i2_3_lut_rep_286_4_lut.init = 16'h6996;
    LUT4 i3_4_lut_adj_302 (.A(block_new_127__N_1901[28]), .B(n33789), .C(n33778), 
         .D(block_new_127__N_1901[12]), .Z(n11918)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i3_4_lut_adj_302.init = 16'h6996;
    LUT4 i27851_2_lut (.A(n6362[3]), .B(n6362[2]), .Z(n30146)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(409[27:47])
    defparam i27851_2_lut.init = 16'heeee;
    LUT4 i4_4_lut_adj_303 (.A(n33584), .B(n33765), .C(block_new_127__N_1901[25]), 
         .D(n33826), .Z(n10_adj_7867)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i4_4_lut_adj_303.init = 16'h6996;
    LUT4 i3_3_lut_4_lut_adj_304 (.A(block_new_127__N_1901[71]), .B(n33803), 
         .C(block_new_127__N_1901[78]), .D(n29244), .Z(n8_adj_7701)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i3_3_lut_4_lut_adj_304.init = 16'h6996;
    LUT4 i1_2_lut_3_lut_adj_305 (.A(block_new_127__N_1901[125]), .B(block_new_127__N_1901[127]), 
         .C(n29231), .Z(n4_adj_7826)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_3_lut_adj_305.init = 16'h9696;
    LUT4 i2_2_lut_3_lut_4_lut_adj_306 (.A(block_new_127__N_1901[51]), .B(n33805), 
         .C(n29408), .D(n11890), .Z(n6_adj_7966)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i2_2_lut_3_lut_4_lut_adj_306.init = 16'h6996;
    LUT4 i1_2_lut_3_lut_4_lut_adj_307 (.A(block_new_127__N_1901[101]), .B(block_new_127__N_1901[103]), 
         .C(block_new_127__N_1901[127]), .D(block_new_127__N_1901[125]), 
         .Z(n6_adj_8020)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_3_lut_4_lut_adj_307.init = 16'h6996;
    LUT4 i6_4_lut (.A(block_new_127__N_1901[66]), .B(n12_adj_8024), .C(block_new_127__N_1901[87]), 
         .D(block_new_127__N_1901[88]), .Z(n29146)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i6_4_lut.init = 16'h6996;
    LUT4 i5_4_lut_adj_308 (.A(block_new_127__N_1901[82]), .B(block_new_127__N_1901[72]), 
         .C(n33762), .D(block_new_127__N_1901[71]), .Z(n12_adj_8024)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i5_4_lut_adj_308.init = 16'h6996;
    LUT4 i3_3_lut (.A(n33581), .B(block_new_127__N_1901[112]), .C(block_new_127__N_1901[121]), 
         .Z(n8_adj_7848)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i3_3_lut.init = 16'h9696;
    LUT4 i1_2_lut_3_lut_4_lut_adj_309 (.A(n33808), .B(n33807), .C(block_new_127__N_1901[100]), 
         .D(block_new_127__N_1901[125]), .Z(n4_adj_7959)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_3_lut_4_lut_adj_309.init = 16'h6996;
    LUT4 i4_4_lut_adj_310 (.A(block_new_127__N_1901[34]), .B(n33694), .C(n33810), 
         .D(n33709), .Z(n10_adj_7834)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i4_4_lut_adj_310.init = 16'h6996;
    LUT4 i4_4_lut_adj_311 (.A(block_new_127__N_1901[33]), .B(block_new_127__N_1901[50]), 
         .C(block_new_127__N_1901[57]), .D(block_new_127__N_1901[42]), .Z(n10_adj_7831)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i4_4_lut_adj_311.init = 16'h6996;
    LUT4 i3_4_lut_adj_312 (.A(block_new_127__N_1901[48]), .B(n33676), .C(block_new_127__N_1901[32]), 
         .D(block_new_127__N_1901[58]), .Z(n29390)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i3_4_lut_adj_312.init = 16'h6996;
    LUT4 i3_3_lut_4_lut_adj_313 (.A(block_new_127__N_1901[122]), .B(block_new_127__N_1901[127]), 
         .C(block_new_127__N_1901[107]), .D(n29220), .Z(n8_adj_7889)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i3_3_lut_4_lut_adj_313.init = 16'h6996;
    LUT4 i1_2_lut_3_lut_adj_314 (.A(block_new_127__N_1901[122]), .B(block_new_127__N_1901[127]), 
         .C(block_new_127__N_1901[115]), .Z(n5_adj_7994)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_3_lut_adj_314.init = 16'h9696;
    LUT4 i1_2_lut_4_lut_adj_315 (.A(n33809), .B(block_new_127__N_1901[83]), 
         .C(block_new_127__N_1901[75]), .D(n33821), .Z(n4_adj_7971)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_4_lut_adj_315.init = 16'h6996;
    LUT4 i1_2_lut_4_lut_adj_316 (.A(n33809), .B(block_new_127__N_1901[83]), 
         .C(block_new_127__N_1901[75]), .D(n29172), .Z(n5_adj_7946)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_4_lut_adj_316.init = 16'h6996;
    LUT4 i2_3_lut_rep_410_4_lut (.A(block_new_127__N_1901[122]), .B(block_new_127__N_1901[127]), 
         .C(n33833), .D(n29339), .Z(n33714)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i2_3_lut_rep_410_4_lut.init = 16'h6996;
    LUT4 i3_3_lut_adj_317 (.A(n29146), .B(block_new_127__N_1901[65]), .C(block_new_127__N_1901[73]), 
         .Z(n8_adj_7795)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i3_3_lut_adj_317.init = 16'h9696;
    LUT4 i4_4_lut_adj_318 (.A(n33680), .B(n12074), .C(block_new_127__N_1901[81]), 
         .D(n33803), .Z(n10_adj_7792)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i4_4_lut_adj_318.init = 16'h6996;
    LUT4 i2_2_lut_3_lut_adj_319 (.A(block_new_127__N_1901[106]), .B(block_new_127__N_1901[111]), 
         .C(n29220), .Z(n7_adj_7992)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i2_2_lut_3_lut_adj_319.init = 16'h9696;
    LUT4 i5_4_lut_adj_320 (.A(block_new_127__N_1901[33]), .B(n33813), .C(block_new_127__N_1901[34]), 
         .D(n29393), .Z(n12)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i5_4_lut_adj_320.init = 16'h6996;
    LUT4 i3_4_lut_adj_321 (.A(block_new_127__N_1901[90]), .B(n33669), .C(n33682), 
         .D(n33771), .Z(n29396)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i3_4_lut_adj_321.init = 16'h6996;
    LUT4 i2_3_lut_rep_411_4_lut (.A(block_new_127__N_1901[98]), .B(block_new_127__N_1901[103]), 
         .C(block_new_127__N_1901[102]), .D(n33835), .Z(n33715)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i2_3_lut_rep_411_4_lut.init = 16'h6996;
    LUT4 i4_4_lut_adj_322 (.A(n33819), .B(block_new_127__N_1901[79]), .C(block_new_127__N_1901[65]), 
         .D(n33804), .Z(n10_adj_7759)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i4_4_lut_adj_322.init = 16'h6996;
    LUT4 i4_4_lut_adj_323 (.A(n33780), .B(block_new_127__N_1901[1]), .C(n6345[3]), 
         .D(n33673), .Z(n10_adj_7746)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i4_4_lut_adj_323.init = 16'h6996;
    LUT4 i4_4_lut_adj_324 (.A(n33698), .B(block_new_127__N_1901[46]), .C(n33799), 
         .D(block_new_127__N_1901[61]), .Z(n10_adj_7740)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i4_4_lut_adj_324.init = 16'h6996;
    LUT4 i1_2_lut_3_lut_adj_325 (.A(block_new_127__N_1901[114]), .B(block_new_127__N_1901[119]), 
         .C(block_new_127__N_1901[107]), .Z(n29441)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i1_2_lut_3_lut_adj_325.init = 16'h9696;
    LUT4 i4_4_lut_adj_326 (.A(n33786), .B(n4770[4]), .C(block_new_127__N_1901[46]), 
         .D(n33802), .Z(n10_adj_7736)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(126[14:31])
    defparam i4_4_lut_adj_326.init = 16'h6996;
    LUT4 i4_4_lut_adj_327 (.A(n33776), .B(block_new_127__N_1901[25]), .C(n33750), 
         .D(block_new_127__N_1901[1]), .Z(n10_adj_7711)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i4_4_lut_adj_327.init = 16'h6996;
    LUT4 i1_2_lut_rep_221_3_lut (.A(block_new_127__N_1901[117]), .B(block_new_127__N_1901[124]), 
         .C(n29160), .Z(n33525)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i1_2_lut_rep_221_3_lut.init = 16'h9696;
    LUT4 i4_4_lut_adj_328 (.A(n33765), .B(block_new_127__N_1901[17]), .C(block_new_127__N_1901[24]), 
         .D(block_new_127__N_1901[15]), .Z(n10)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(120[14:31])
    defparam i4_4_lut_adj_328.init = 16'h6996;
    LUT4 i3_4_lut_adj_329 (.A(block_new_127__N_1901[38]), .B(block_new_127__N_1901[34]), 
         .C(block_new_127__N_1901[49]), .D(block_new_127__N_1901[42]), .Z(n28987)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i3_4_lut_adj_329.init = 16'h6996;
    LUT4 i2_2_lut_3_lut_adj_330 (.A(block_new_127__N_1901[123]), .B(block_new_127__N_1901[127]), 
         .C(block_new_127__N_1901[116]), .Z(n7_adj_7996)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/suhail/downloads/aes-master/aes-master/src/rtl/aes_decipher_block.v(84[13:53])
    defparam i2_2_lut_3_lut_adj_330.init = 16'h9696;
    PFUMX mux_625_i120 (.BLUT(n2_adj_8016), .ALUT(n4540[119]), .C0(n30026), 
          .Z(n3899[119]));
    PFUMX mux_625_i115 (.BLUT(n2_adj_8015), .ALUT(n4540[114]), .C0(n30026), 
          .Z(n3899[114]));
    PFUMX mux_625_i88 (.BLUT(n2_adj_8014), .ALUT(n4540[87]), .C0(n30026), 
          .Z(n3899[87]));
    PFUMX mux_625_i73 (.BLUT(n2_adj_8013), .ALUT(n4540[72]), .C0(n30026), 
          .Z(n3899[72]));
    PFUMX mux_625_i66 (.BLUT(n2_adj_8011), .ALUT(n4540[65]), .C0(n30026), 
          .Z(n3899[65]));
    PFUMX mux_625_i59 (.BLUT(n2_adj_8009), .ALUT(n4540[58]), .C0(n30026), 
          .Z(n3899[58]));
    PFUMX mux_625_i56 (.BLUT(n2_adj_8007), .ALUT(n4540[55]), .C0(n30026), 
          .Z(n3899[55]));
    PFUMX mux_625_i49 (.BLUT(n2_adj_8006), .ALUT(n4540[48]), .C0(n30026), 
          .Z(n3899[48]));
    PFUMX mux_625_i24 (.BLUT(n2_adj_8004), .ALUT(n4540[23]), .C0(n30026), 
          .Z(n3899[23]));
    PFUMX mux_625_i8 (.BLUT(n2_adj_8019), .ALUT(n4540[7]), .C0(n30026), 
          .Z(n3899[7]));
    
endmodule

/******************************************************************************
Copyright 2017 Gnarly Grey LLC

Permission is hereby granted, free of charge, to any person obtaining a copy
of this software and associated documentation files (the "Software"), to deal
in the Software without restriction, including without limitation the rights
to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
copies of the Software, and to permit persons to whom the Software is
furnished to do so, subject to the following conditions:

The above copyright notice and this permission notice shall be included in all
copies or substantial portions of the Software.

THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
SOFTWARE.
******************************************************************************/

module ebr_bm_mem (
  input           clk,
  input  [4:0]    bm_no,
  input  [8:0]    addr,
  output [7:0]    data
  );

  reg    [23:0]   read_en;
  reg    [7:0]    data_reg;
  wire   [7:0]    data_int[23:0];
  
  assign          data = data_reg;
  
  always @ (posedge clk)
    begin
      read_en <= 24'h000000;
      case (bm_no)
        5'd0    : read_en[0]  <= 1'b1;
        5'd1    : read_en[1]  <= 1'b1;
        5'd2    : read_en[2]  <= 1'b1;
        5'd3    : read_en[3]  <= 1'b1;
        5'd4    : read_en[4]  <= 1'b1;
        5'd5    : read_en[5]  <= 1'b1;
        5'd6    : read_en[6]  <= 1'b1;
        5'd7    : read_en[7]  <= 1'b1;
        5'd8    : read_en[8]  <= 1'b1;
        5'd9    : read_en[9]  <= 1'b1;
        5'd10   : read_en[10] <= 1'b1;
        5'd11   : read_en[11] <= 1'b1;
        5'd12   : read_en[12] <= 1'b1;
        5'd13   : read_en[13] <= 1'b1;
        5'd14   : read_en[14] <= 1'b1;
        5'd15   : read_en[15] <= 1'b1;
        5'd16   : read_en[16] <= 1'b1;
        5'd17   : read_en[17] <= 1'b1;
        5'd18   : read_en[18] <= 1'b1;
        5'd19   : read_en[19] <= 1'b1;
        5'd20   : read_en[20] <= 1'b1;
        5'd21   : read_en[21] <= 1'b1;
        5'd22   : read_en[22] <= 1'b1;
        5'd23   : read_en[23] <= 1'b1;        
        default : read_en[0]  <= 1'b1;
      endcase
    end
  
  always @ (*)
    begin
      case (bm_no)
        5'd0    : data_reg <= data_int[0] ;
        5'd1    : data_reg <= data_int[1] ;
        5'd2    : data_reg <= data_int[2] ;
        5'd3    : data_reg <= data_int[3] ;
        5'd4    : data_reg <= data_int[4] ;
        5'd5    : data_reg <= data_int[5] ;
        5'd6    : data_reg <= data_int[6] ;
        5'd7    : data_reg <= data_int[7] ;
        5'd8    : data_reg <= data_int[8] ;
        5'd9    : data_reg <= data_int[9] ;
        5'd10   : data_reg <= data_int[10];
        5'd11   : data_reg <= data_int[11];
        5'd12   : data_reg <= data_int[12];
        5'd13   : data_reg <= data_int[13];
        5'd14   : data_reg <= data_int[14];
        5'd15   : data_reg <= data_int[15];
        5'd16   : data_reg <= data_int[16];
        5'd17   : data_reg <= data_int[17];
        5'd18   : data_reg <= data_int[18];
        5'd19   : data_reg <= data_int[19];
        5'd20   : data_reg <= data_int[20];
        5'd21   : data_reg <= data_int[21];
        5'd22   : data_reg <= data_int[22];
        5'd23   : data_reg <= data_int[23];        
        default : data_reg <= data_int[0] ;      
      endcase
    end    
  
  SB_RAM512x8 bm0 (
    .RDATA (data_int[0]),
    .RADDR (addr),
    .RCLK  (clk),
    .RCLKE (read_en[0]),
    .RE    (read_en[0]),
    .WADDR (9'h000),
    .WCLK  (1'b0),
    .WCLKE (1'b0),
    .WDATA (8'h00),
    .WE    (1'b0)
  );  
  defparam bm0.INIT_0 = 256'h00003e007e0000000000fcf71f0000000000f0ff07000000000080ff01000000;
  defparam bm0.INIT_1 = 256'h00e001008007000000c00300c003000000800700e001000000001f00f8000000;
  defparam bm0.INIT_2 = 256'h00380000001e000000780000000e000000700000000e000000f0000000070000;
  defparam bm0.INIT_3 = 256'h801f000000001f00001c000000f80f00001c000000fc03000038000000fc0000;
  defparam bm0.INIT_4 = 256'h3c1c00000000801f781c00000000f007f01d00000000f803e01f000000007c00;
  defparam bm0.INIT_5 = 256'h07380000000000700f380000000000700e1c0000000000381c1c00000000003e;
  defparam bm0.INIT_6 = 256'h07e00100000000e007f00000000000e007700000000000e007780000000000e0;
  defparam bm0.INIT_7 = 256'h0e003e00000000e007000f00000000e007800700000000e007c00300000000e0;
  defparam bm0.INIT_8 = 256'hf80000000000001e3c00c00f0000003c1c00f00f000000780e00fc0300000070;
  defparam bm0.INIT_9 = 256'h00f8ffffffff1f0080ffffffffffff01c0ffffffffffff07f00700000000c00f;
  defparam bm0.INIT_A = 256'h00f81d0000b81f0000f81d0000b81f00000018000018000000003800001c0000;
  defparam bm0.INIT_B = 256'h00003800001c000000003800001c000000001c000038000000f81d0000b81f00;
  defparam bm0.INIT_C = 256'h0080e0018007010000c0f30000cf030000c0730000ce030000003b0000dc0000;
  defparam bm0.INIT_D = 256'h00003cfc3f3c0000000038ffff1c00000000900ff00900000000c003c0030000;
  defparam bm0.INIT_E = 256'h00000087e100000000000687e160000000000e066070000000001ef00f780000;
  defparam bm0.INIT_F = 256'h00000080010000000000008001000000000000800100000000000083c1000000;

  SB_RAM512x8 bm1 (
    .RDATA (data_int[1]),
    .RADDR (addr),
    .RCLK  (clk),
    .RCLKE (read_en[1]),
    .RE    (read_en[1]),
    .WADDR (9'h000),
    .WCLK  (1'b0),
    .WCLKE (1'b0),
    .WDATA (8'h00),
    .WE    (1'b0)
  );  
  defparam bm1.INIT_0 = 256'h0000b807007007000000f80300f007000000f00300f007000000f00100e00300;
  defparam bm1.INIT_1 = 256'h00f8ffffffffff07000038070070070000003807007007000000380700700700;
  defparam bm1.INIT_2 = 256'h001c00000000001e001c00000000001e00fcffffffffff1f00fcffffffffff0f;
  defparam bm1.INIT_3 = 256'h001c00000000001e001c00000000001e001c00000000001e001c00000000001e;
  defparam bm1.INIT_4 = 256'h00fcffffffff1f1e00fcffffffff3f1e00fcffffffff3f1e001c00000000001e;
  defparam bm1.INIT_5 = 256'h001cfc877ff80f1e001c00000000001e001c00000000001e001c00000000001e;
  defparam bm1.INIT_6 = 256'h001cfcc7fff80f1e001c1cc7e3380e1e001cfcc7fff80f1e001cfcc7fff80f1e;
  defparam bm1.INIT_7 = 256'h001c00000000001e001c00000000001e001cfc877ff80f1e001cfcc7fff80f1e;
  defparam bm1.INIT_8 = 256'h0000fcc7fff80f1e000cfc877ff80f1e001c00000000001e001c00000000001e;
  defparam bm1.INIT_9 = 256'h00feffc7fff80f1e00f8ffc7fff80f1e00e03fc7e3380e1e0000fcc7fff80f1e;
  defparam bm1.INIT_A = 256'he001001e0000001ec003001f0000001e800f800f0000001e001fe0877ff80f1e;
  defparam bm1.INIT_B = 256'h708003f0e3380e1e708003f8fff80f1ef08003b8fff80f1ee081033c7ff0071e;
  defparam bm1.INIT_C = 256'h708007f07ff80f1e788003f0fff80f1e708003f0fff80f1e708003f0e3380e1e;
  defparam bm1.INIT_D = 256'hf00018f8ffffff1f70001c780000001e70001e700000001e70000f700000001e;
  defparam bm1.INIT_E = 256'h800f800f00000000c003001f00000000e00100feffffff0fe00100fcffffff1f;
  defparam bm1.INIT_F = 256'h00e03f000000000000f8ff000000000000feff0300000000001fe00700000000;

  SB_RAM512x8 bm2 (
    .RDATA (data_int[2]),
    .RADDR (addr),
    .RCLK  (clk),
    .RCLKE (read_en[2]),
    .RE    (read_en[2]),
    .WADDR (9'h000),
    .WCLK  (1'b0),
    .WCLKE (1'b0),
    .WDATA (8'h00),
    .WE    (1'b0)
  );  
  defparam bm2.INIT_0 = 256'hfffffffffffffffffffffffffffffffffeffffffffffff7ffcffffffffffff3f;
  defparam bm2.INIT_1 = 256'h0f000000000000f00f000000000000f00f000000000000f00f000000000000f0;
  defparam bm2.INIT_2 = 256'h0f809f9f03fffcf00ffe1f8ff7fff8f00ffe1f8ffffff0f00f780c06fb6760f0;
  defparam bm2.INIT_3 = 256'h0f1ff8fbe1fff7f00ffef9fff9fffff00ff8bbdff9fffef00fc0bfdf03fffef0;
  defparam bm2.INIT_4 = 256'h0ffce070f8e7e0f00ffef1f0f8fff1f00ffff1f900fff1f00f0ff0f900fff3f0;
  defparam bm2.INIT_5 = 256'h0f000000000000f00f000000000000f00f000000000000f00f000000000000f0;
  defparam bm2.INIT_6 = 256'hcffffffffffffff38ffffffffffffff18ffffffffffffff10f000000000000f0;
  defparam bm2.INIT_7 = 256'h0f000000000000f00f000000000000f00f000000000000f08ffffffffffffff1;
  defparam bm2.INIT_8 = 256'h8ffffffffffffff10ffffffffffffff00f000000000000f00f000000000000f0;
  defparam bm2.INIT_9 = 256'h0f000000000000f00ffeffffffff7ff08ffffffffffffff1cffffffffffffff3;
  defparam bm2.INIT_A = 256'h0ffffffffffffff00f000000000000f00f000000000000f00f000000000000f0;
  defparam bm2.INIT_B = 256'h0ffffffffffffff08ffffffffffffff1cffffffffffffff38ffffffffffffff1;
  defparam bm2.INIT_C = 256'hffffff03000000f00f000000000000f00f000000000000f00f000000000000f0;
  defparam bm2.INIT_D = 256'hf83f80c7fffffff1feffffc7fffffff3feffffc7fffffff1ffffff07000000f0;
  defparam bm2.INIT_E = 256'h00f0ff07000000f000fc9f07000000f000ff8707000000f0e0ff8087fffffff1;
  defparam bm2.INIT_F = 256'h0000c0ffffffff3f0000f0ffffffff7f0000feffffffffff0080ffffffffffff;

  SB_RAM512x8 bm3 (
    .RDATA (data_int[3]),
    .RADDR (addr),
    .RCLK  (clk),
    .RCLKE (read_en[3]),
    .RE    (read_en[3]),
    .WADDR (9'h000),
    .WCLK  (1'b0),
    .WCLKE (1'b0),
    .WDATA (8'h00),
    .WE    (1'b0)
  );  
  defparam bm3.INIT_0 = 256'h00c003c003c0030000c003c003c0030000c003c003c0030000c003c003c00300;
  defparam bm3.INIT_1 = 256'hfeffffffffffff7ffcffffffffffff3f00c003c003c0030000c003c003c00300;
  defparam bm3.INIT_2 = 256'h0fc003c003c003f01fc003c003c003f8ffffffffffffffffffffffffffffffff;
  defparam bm3.INIT_3 = 256'h0fc003c003c003f00fc003c003c003f00fc003c003c003f00fc003c003c003f0;
  defparam bm3.INIT_4 = 256'h0f000000000000f00f000000000000f00f000000000000f00f000000000000f0;
  defparam bm3.INIT_5 = 256'h0f000000000000f00f000000000000f00f000000000000f00f000000000000f0;
  defparam bm3.INIT_6 = 256'h0fc03ff00ffc03f00fc03ff00ffc03f00fc03ff00ffc03f00fc03ff00ffc03f0;
  defparam bm3.INIT_7 = 256'h0f000000000000f00f000000000000f00fc03ff00ffc03f00fc03ff00ffc03f0;
  defparam bm3.INIT_8 = 256'h0fc03ff00ffc03f00fc03ff00ffc03f00f000000000000f00f000000000000f0;
  defparam bm3.INIT_9 = 256'h0fc03ff00ffc03f00fc03ff00ffc03f00fc03ff00ffc03f00fc03ff00ffc03f0;
  defparam bm3.INIT_A = 256'h0f000000000000f00f000000000000f00f000000000000f00f000000000000f0;
  defparam bm3.INIT_B = 256'h0fc03ff00ffc03f00fc03ff00ffc03f00fc03ff00ffc03f00fc03ff00ffc03f0;
  defparam bm3.INIT_C = 256'h0f000000000000f00f000000000000f00fc03ff00ffc03f00fc03ff00ffc03f0;
  defparam bm3.INIT_D = 256'h0f000000000000f00f000000000000f00f000000000000f00f000000000000f0;
  defparam bm3.INIT_E = 256'h1f000000000000f80f000000000000f00f000000000000f00f000000000000f0;
  defparam bm3.INIT_F = 256'hfcffffffffffff3ffeffffffffffff7fffffffffffffffffffffffffffffffff;

  SB_RAM512x8 bm4 (
    .RDATA (data_int[4]),
    .RADDR (addr),
    .RCLK  (clk),
    .RCLKE (read_en[4]),
    .RE    (read_en[4]),
    .WADDR (9'h000),
    .WCLK  (1'b0),
    .WCLKE (1'b0),
    .WDATA (8'h00),
    .WE    (1'b0)
  );  
  defparam bm4.INIT_0 = 256'h80f0ffffffff0f010070000000000e0000f0ffffffff0f0000f0ffffffff0f00;
  defparam bm4.INIT_1 = 256'h0e600000000006701e78000000001e78fc7f00000000fe3ff0ffffffffffff0f;
  defparam bm4.INIT_2 = 256'h3be00000000007dc77f8000000001feef7ff00000000ffefe77f00000000ffe7;
  defparam bm4.INIT_3 = 256'h33c00000000003cc3bc00000000003dc3be00000000007dc3be00000000007dc;
  defparam bm4.INIT_4 = 256'h77c00100008003ee77c00100008003ee77c00100008003ee77c00100008003ee;
  defparam bm4.INIT_5 = 256'hdc81030000d8813bce81030000f88173ee80030000f80177e680010000b00167;
  defparam bm4.INIT_6 = 256'h701e0e00007e780e780f070000fcf01eb807070000fce01d9c03030000dcc039;
  defparam bm4.INIT_7 = 256'h80cf3f0080fff30180f31f0000fecf01c0f90c0000379f03e03c0e00007e3c07;
  defparam bm4.INIT_8 = 256'h00c0ff0180ff030000f0ff0000ff0f0000fc7000800f3f00003e3c00c03d7c00;
  defparam bm4.INIT_9 = 256'h003e001c38000000000c000ff000000000008007e00100030000fe03c07f0003;
  defparam bm4.INIT_A = 256'h000c00fc3f700000000c00fc3f700000003f00f81f700000003f00381c000000;
  defparam bm4.INIT_B = 256'h008003f81f000000000000fc3f0000000000000e700000000000000e70000000;
  defparam bm4.INIT_C = 256'h000080ffff017c00000000381c007c00000003381c007c00008003381c001800;
  defparam bm4.INIT_D = 256'h0000c001800300000000c001800300000000c0ffff0300000000c0ffff033800;
  defparam bm4.INIT_E = 256'h00000e000070000000000e00007000000000feffff7f00000000feffff7f0000;
  defparam bm4.INIT_F = 256'h0000feffff7f00000000feffff7f000000000e000070000000000e0000700000;

  SB_RAM512x8 bm5 (
    .RDATA (data_int[5]),
    .RADDR (addr),
    .RCLK  (clk),
    .RCLKE (read_en[5]),
    .RE    (read_en[5]),
    .WADDR (9'h000),
    .WCLK  (1'b0),
    .WCLKE (1'b0),
    .WDATA (8'h00),
    .WE    (1'b0)
  );  
  defparam bm5.INIT_0 = 256'h000000c0c707000000000080ff03000000000000ff01000000000000fe000000;
  defparam bm5.INIT_1 = 256'h000000e0010f0000000000e0010f0000000000e0010f0000000000c083070000;
  defparam bm5.INIT_2 = 256'h000000e0010f000000e0ffe1010f000000e0ffe1010f000000e0ffe1010f0000;
  defparam bm5.INIT_3 = 256'h0000fce1010f00000000fce1010f0000000000e0010f0000000000e0010f0000;
  defparam bm5.INIT_4 = 256'h000000e0010f0000000000e0010f0000000000e0010f00000000fce1010f0000;
  defparam bm5.INIT_5 = 256'h000000e0010f000000e0ffe1010f000000e0ffe1010f000000e0ffe1010f0000;
  defparam bm5.INIT_6 = 256'h0000fce17d0f00000000fce17d0f0000000000e07d0f0000000000e0390f0000;
  defparam bm5.INIT_7 = 256'h000000e07d0f0000000000e07d0f0000000000e07d0f00000000fce17d0f0000;
  defparam bm5.INIT_8 = 256'h000000e07d0f000000e0ffe17d0f000000e0ffe17d0f000000e0ffe17d0f0000;
  defparam bm5.INIT_9 = 256'h000000f87d3f0000000000e07d0f0000000000e07d0f0000000000e07d0f0000;
  defparam bm5.INIT_A = 256'h000000cfdfe701000000001efff100000000003e7cf80000000000fc7c7e0000;
  defparam bm5.INIT_B = 256'h000080f3ff980300000080f33fdc0300000080e71fcc0300000000e70fce0100;
  defparam bm5.INIT_C = 256'h0000c0f3ff9f07000000c0fbffb907000000c0fbffb807000000c0f3ff980300;
  defparam bm5.INIT_D = 256'h000080e7ffcf0300000080e7ffcf0300000080f3ffdf0300000080f3ff9f0300;
  defparam bm5.INIT_E = 256'h0000007c007e00000000003efef800000000009ffff30100000000cfffe70100;
  defparam bm5.INIT_F = 256'h00000000ff010000000000c0ff070000000000f0ff1f0000000000f8c73f0000;  
  
  SB_RAM512x8 bm6 (
    .RDATA (data_int[6]),
    .RADDR (addr),
    .RCLK  (clk),
    .RCLKE (read_en[6]),
    .RE    (read_en[6]),
    .WADDR (9'h000),
    .WCLK  (1'b0),
    .WCLKE (1'b0),
    .WDATA (8'h00),
    .WE    (1'b0)
  );  
  defparam bm6.INIT_0 = 256'h0000800ff8000000000080ffff000000000000ff7f000000000000fc1f000000;
  defparam bm6.INIT_1 = 256'h0000c0f3ef0100000000c003e00100000000c003e001000000008007f0010000;
  defparam bm6.INIT_2 = 256'h0000f00ff00f00000000e0ffff0700000000c0ffff0100000000c0ffff010000;
  defparam bm6.INIT_3 = 256'h00000f0000f8000000003f0000fc000000007e00007e00000000fc01803f0000;
  defparam bm6.INIT_4 = 256'h00e00100f0c1070000c00300f8c0030000c0070078e003000080070000f00100;
  defparam bm6.INIT_5 = 256'h00f0000080070f0000f00000c0070f0000f00000c0830f0000e00100e0810700;
  defparam bm6.INIT_6 = 256'h00780000000f1e0000780000000f0e0000700000000f0f000070000080070f00;
  defparam bm6.INIT_7 = 256'h00780000000e1e0000780000000e1e0000780000000f1e0000780000000f1e00;
  defparam bm6.INIT_8 = 256'h00380000001e1c0000380000001e1e0000380000000e1e0000780000000e1e00;
  defparam bm6.INIT_9 = 256'h003c0000001e3c00003c0000001e3c00003c0000001e3c00003c0000001e3c00;
  defparam bm6.INIT_A = 256'h001e000000007800001e0000001c7800001e0000001c7800001c0000001e3c00;
  defparam bm6.INIT_B = 256'h800700000078f001000f00000078f000000f00000030f000000f000000007800;
  defparam bm6.INIT_C = 256'hc00300000000c003c00300000000c003800300000000e001800700000030e001;
  defparam bm6.INIT_D = 256'h80ffffffffffff01c0ffffffffffff03c0ffffffffffff03c001000000008003;
  defparam bm6.INIT_E = 256'h0000001ff80000000000000ff00000000000000ff000000000ffffffffffff00;
  defparam bm6.INIT_F = 256'h000000f00f000000000000f81f000000000000fc3f0000000000007e7f000000;

  SB_RAM512x8 bm7 (
    .RDATA (data_int[7]),
    .RADDR (addr),
    .RCLK  (clk),
    .RCLKE (read_en[7]),
    .RE    (read_en[7]),
    .WADDR (9'h000),
    .WCLK  (1'b0),
    .WCLKE (1'b0),
    .WDATA (8'h00),
    .WE    (1'b0)
  );  
  defparam bm7.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam bm7.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam bm7.INIT_2 = 256'hfffffffffffffffffeffffffffffff7ffcffffffffffff1f0000000000000000;
  defparam bm7.INIT_3 = 256'h3f000000000000fc1f000000000000f00f000000000000f0ffffffffffffffff;
  defparam bm7.INIT_4 = 256'he70700000000e0e7f7030000000080ffff000000000000ff7f000000000000fe;
  defparam bm7.INIT_5 = 256'h07fc000000003fe0077e000000007ee0073f00000000f8e1c70f00000000f0e3;
  defparam bm7.INIT_6 = 256'h07801f0000f801e007c00f0000f003e007e0070000c00fe007f8010000801fe0;
  defparam bm7.INIT_7 = 256'h0700f007c00f00e00700f801801f00e00700fc00003f00e007007e0000fc00e0;
  defparam bm7.INIT_8 = 256'h0700f0ffff0f00e00700e03ffc0700e00700801ff80100e00700c00fe00700e0;
  defparam bm7.INIT_9 = 256'h07801f0000f801e007003fc003fc00e00700fcf00f3f00e00700f8f99f1f00e0;
  defparam bm7.INIT_A = 256'h07fc000000003fe007f8010000801fe007f0030000e00fe007c00f0000f003e0;
  defparam bm7.INIT_B = 256'he70700000000e0e7c70f00000000f0e3871f00000000f8e1077e000000007ee0;
  defparam bm7.INIT_C = 256'h3f000000000000fc7f000000000000feff000000000000ffff0100000000c0ff;
  defparam bm7.INIT_D = 256'h0000000000000000f8ffffffffffff1ffeffffffffffff7fffffffffffffffff;
  defparam bm7.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam bm7.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

  SB_RAM512x8 bm8 (
    .RDATA (data_int[8]),
    .RADDR (addr),
    .RCLK  (clk),
    .RCLKE (read_en[8]),
    .RE    (read_en[8]),
    .WADDR (9'h000),
    .WCLK  (1'b0),
    .WCLKE (1'b0),
    .WDATA (8'h00),
    .WE    (1'b0)
  );  
  defparam bm8.INIT_0 = 256'h0000008001000000000000800100000000000080010000000000008001000000;
  defparam bm8.INIT_1 = 256'h00007080010e000000007080010e000000000080010000000000008001000000;
  defparam bm8.INIT_2 = 256'h001c40f00f023800000ec000000370000006e080010760000000e08001070000;
  defparam bm8.INIT_3 = 256'h00c0f900009f030000e0f007e00f07000070c0ffff030e00003800ffff001c00;
  defparam bm8.INIT_4 = 256'h0080070000e0010000000f0000f0000000001e000078000000807c00003e0100;
  defparam bm8.INIT_5 = 256'h00e700000000e700c0ef01000080f703c0c301000080c303c0c0030000c00303;
  defparam bm8.INIT_6 = 256'h0030000000000c000070000000000e000070000000000e000070000000000e00;
  defparam bm8.INIT_7 = 256'hff3b00000000dcff0038000000001c000038000000001c000038000000001c00;
  defparam bm8.INIT_8 = 256'h0038000000001c000038000000001c000038000000001c00ff3b00000000dcff;
  defparam bm8.INIT_9 = 256'h0070000000000e000070000000000e000070000000000e000030000000000c00;
  defparam bm8.INIT_A = 256'hc0c0030000c00303c0c301000080c303c0ef01000080f70300e700000000e700;
  defparam bm8.INIT_B = 256'h00807c00003e010000001e000078000000000f0000f000000080070000e00100;
  defparam bm8.INIT_C = 256'h003800ffff001c000070c0ffff030e0000e0f007e00f070000c0f900009f0300;
  defparam bm8.INIT_D = 256'h0000e080010700000006e08001076000000ec00000037000001c40f00f023800;
  defparam bm8.INIT_E = 256'h0000008001000000000000800100000000007080010e000000007080010e0000;
  defparam bm8.INIT_F = 256'h0000008001000000000000800100000000000080010000000000008001000000;

  SB_RAM512x8 bm9 (
    .RDATA (data_int[9]),
    .RADDR (addr),
    .RCLK  (clk),
    .RCLKE (read_en[9]),
    .RE    (read_en[9]),
    .WADDR (9'h000),
    .WCLK  (1'b0),
    .WCLKE (1'b0),
    .WDATA (8'h00),
    .WE    (1'b0)
  );  
  defparam bm9.INIT_0 = 256'h0080f7f0807f000000001c70ff1f000000001cf0ff03000000001cf07f000000;
  defparam bm9.INIT_1 = 256'h00001c001e001f0000001c000f800f000000ffc007e003000080f7e003fc0100;
  defparam bm9.INIT_2 = 256'h000000007000e001000000007000f0000000000078007800000018003c003c00;
  defparam bm9.INIT_3 = 256'h001cc01fc001000f001c0007c001000700000006e000800300000000e000c003;
  defparam bm9.INIT_4 = 256'h80ff00078001003880f700078001001c80ffc01fc001001c001cc01dc001000e;
  defparam bm9.INIT_5 = 256'h0000000080010070001c000080010070001c000080030070001c000080030038;
  defparam bm9.INIT_6 = 256'h00000000e00000e000000000c00100e000000000c00100e000000000c0010070;
  defparam bm9.INIT_7 = 256'h3f000000780000e03f000000700000e01f000000e00000e000000000e00000e0;
  defparam bm9.INIT_8 = 256'hc7030080070000e0e70100000e0000e0f70000001c0000e073000000380000e0;
  defparam bm9.INIT_9 = 256'h0ef8ff3f0000006007fc03ff000000e0073f00f0010000e0870f00c0030000e0;
  defparam bm9.INIT_A = 256'h1c000000000000380c000000000000300e000000000000700ec0ff0f00000070;
  defparam bm9.INIT_B = 256'h700000000000000e380000000000001c380000000000001c1c00000000000038;
  defparam bm9.INIT_C = 256'hc00300000000c003e001000000008007e000000000000007f00000000000000f;
  defparam bm9.INIT_D = 256'h003c000000003c00001e000000007800000f00000000f000800700000000e001;
  defparam bm9.INIT_E = 256'h00801f0000f8010000c0070000e0070000f0010000800f0000f8000000001e00;
  defparam bm9.INIT_F = 256'h000000fe7f0000000000e0ffff0700000000f8ffff1f00000000fe01007f0000;

  SB_RAM512x8 bm10 (
    .RDATA (data_int[10]),
    .RADDR (addr),
    .RCLK  (clk),
    .RCLKE (read_en[10]),
    .RE    (read_en[10]),
    .WADDR (9'h000),
    .WCLK  (1'b0),
    .WCLKE (1'b0),
    .WDATA (8'h00),
    .WE    (1'b0)
  );  
  defparam bm10.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam bm10.INIT_1 = 256'h00000000001c000000000000001c000000000000000000000000000000000000;
  defparam bm10.INIT_2 = 256'h00000020781c070200000000381c0e0000000000301c060000000000001c0000;
  defparam bm10.INIT_3 = 256'h000000c0f1ffe701000000e0e1ffc103000000f0007f80070000007030000707;
  defparam bm10.INIT_4 = 256'h0000e0ff0700781e0000003e0f003c00000000003e001e0000000080fc80cf00;
  defparam bm10.INIT_5 = 256'h00800f00f000c00100003f007c00e0000000fc803f00e00c0000f8ff0f00f01e;
  defparam bm10.INIT_6 = 256'h00f00000000fc0fd00e001008007c0fd00c00100c003c0f900c00300e001c001;
  defparam bm10.INIT_7 = 256'h0038000000fce10000380000001cc00100380000000ec00100700000000ec001;
  defparam bm10.INIT_8 = 256'he01f00000000fc00c01f000000007e1c001e000000c87f1e001c000000f8e71e;
  defparam bm10.INIT_9 = 256'h0e1c00000000003c1c1c00000000001e7c1c00000000f00ff81c00000000f807;
  defparam bm10.INIT_A = 256'h07700000000000e007380000000000e007380000000000700e18000000000078;
  defparam bm10.INIT_B = 256'h07c00300000000e007e00100000000c003e00000000000e007700000000000e0;
  defparam bm10.INIT_C = 256'h1e00f80f000000700e007e00000000f007001f00000000e007800700000000e0;
  defparam bm10.INIT_D = 256'he0ffffffffffff0ff80000000000001f7800000f0000003c1c00e00f00000038;
  defparam bm10.INIT_E = 256'h0000000000000000000000000000000000ffffffffffff00c0ffffffffffff03;
  defparam bm10.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

  SB_RAM512x8 bm11 (
    .RDATA (data_int[11]),
    .RADDR (addr),
    .RCLK  (clk),
    .RCLKE (read_en[11]),
    .RE    (read_en[11]),
    .WADDR (9'h000),
    .WCLK  (1'b0),
    .WCLKE (1'b0),
    .WDATA (8'h00),
    .WE    (1'b0)
  );  
  defparam bm11.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam bm11.INIT_1 = 256'h000000001cfc0f00000000000cf8010000000000000000000000000000000000;
  defparam bm11.INIT_2 = 256'h000000001cf0c003000000003f78f00100000000733cfc00000000007ffc3f00;
  defparam bm11.INIT_3 = 256'h00000000c081011c00000000c0c1011e0000000000c0010f000000000ce08007;
  defparam bm11.INIT_4 = 256'h0000e0ffc38103700000003ef0870370000000007087033800000000f0870338;
  defparam bm11.INIT_5 = 256'h00800f00f0c101e000003f007cc001e00000fc803fc003e00000f8ffdf8103e0;
  defparam bm11.INIT_6 = 256'h00f00000003f00e000e00100807f00c000c00100c0f300e000c00300e0e100e0;
  defparam bm11.INIT_7 = 256'h0038000000fc016000380000001c00e000380000000e00e000700000001e00e0;
  defparam bm11.INIT_8 = 256'he01f00000000fc3dc01f000000001e38001e000000c80f70001c000000f80770;
  defparam bm11.INIT_9 = 256'h0e1c00000000003c1c1c00000000001e7c1c00000000f00ff81c00000000f81f;
  defparam bm11.INIT_A = 256'h07700000000000e007380000000000e007380000000000700e18000000000078;
  defparam bm11.INIT_B = 256'h07c00300000000e007e00100000000c003e00000000000e007700000000000e0;
  defparam bm11.INIT_C = 256'h1e00f80f000000700e007e00000000f007001f00000000e007800700000000e0;
  defparam bm11.INIT_D = 256'he0ffffffffffff0ff80000000000001f7800000f0000003c1c00e00f00000038;
  defparam bm11.INIT_E = 256'h0000000000000000000000000000000000ffffffffffff00c0ffffffffffff03;
  defparam bm11.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  
  SB_RAM512x8 bm12 (
    .RDATA (data_int[12]),
    .RADDR (addr),
    .RCLK  (clk),
    .RCLKE (read_en[12]),
    .RE    (read_en[12]),
    .WADDR (9'h000),
    .WCLK  (1'b0),
    .WCLKE (1'b0),
    .WDATA (8'h00),
    .WE    (1'b0)
  );  
  defparam bm12.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam bm12.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam bm12.INIT_2 = 256'h00000080ff3f000000000000ff0f000000000000f80300000000000000000000;
  defparam bm12.INIT_3 = 256'h0000007f00c001000000007000e00100000000e001f00000000000e0077c0000;
  defparam bm12.INIT_4 = 256'h00003f00fc00ff000000fc803f007f000000f8ff0f801f000000e0ff07800300;
  defparam bm12.INIT_5 = 256'h00e000008007003c00e00100c003801f00c00300c001c00f00800f00f000e001;
  defparam bm12.INIT_6 = 256'h00380000001c00e000380000000e00e000700000000e00f000f0000000070078;
  defparam bm12.INIT_7 = 256'hc01f000000001ee0001f000000880fe0001c000000f807e00018000000fc03e0;
  defparam bm12.INIT_8 = 256'h1c1c00000000001e3c1c00000000e03ff81c00000000f87fe01f00000000fcf1;
  defparam bm12.INIT_9 = 256'h07380000000000e007380000000000700e180000000000780e1c00000000003c;
  defparam bm12.INIT_A = 256'h07e00100000000c007e00000000000e007700000000000e007700000000000e0;
  defparam bm12.INIT_B = 256'h0e00fe00000000f007001f00000000e007800700000000e007c00300000000e0;
  defparam bm12.INIT_C = 256'hf00100000000001f7800000f0000003c3c00e00f000000381e00f80f00000070;
  defparam bm12.INIT_D = 256'h000000000000000000feffffffffff0080ffffffffffff03e0ffffffffffff0f;
  defparam bm12.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam bm12.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

  SB_RAM512x8 bm13 (
    .RDATA (data_int[13]),
    .RADDR (addr),
    .RCLK  (clk),
    .RCLKE (read_en[13]),
    .RE    (read_en[13]),
    .WADDR (9'h000),
    .WCLK  (1'b0),
    .WCLKE (1'b0),
    .WDATA (8'h00),
    .WE    (1'b0)
  );  
  defparam bm13.INIT_0 = 256'h00000080ff3f000000000000ff0f000000000000f80300000000000000000000;
  defparam bm13.INIT_1 = 256'h0000007f00c001000000007000e00100000000e001f00000000000e0077c0000;
  defparam bm13.INIT_2 = 256'h00003f007c00ff000000fc803f007f000000f8ff0f800f000000e0ff07800300;
  defparam bm13.INIT_3 = 256'h00e000008007003c00e00100c003801f00c00300c001c00f00800f00f000f001;
  defparam bm13.INIT_4 = 256'h00380000001c00e000380000000e00e000700000000e00f000f0000000070078;
  defparam bm13.INIT_5 = 256'hc01f000000001ee0001f000000880fe0001c000000f807e00018000000fc03e0;
  defparam bm13.INIT_6 = 256'h1c1c00000000001e7c1c00000000e03ff81c00000000f87fe01f00000000fcf1;
  defparam bm13.INIT_7 = 256'h07380000000000e007380000000000700e180000000000780e1c00000000003c;
  defparam bm13.INIT_8 = 256'h07e00100000000c003e00000000000e007700000000000e007700000000000e0;
  defparam bm13.INIT_9 = 256'h0e00fe00000000f007001f00000000e007800700000000e007c00300000000e0;
  defparam bm13.INIT_A = 256'hf00100000000001f7800000f0000003c3c00e00f000000381e00f80f00000070;
  defparam bm13.INIT_B = 256'h000087c3c1e10000009e83c3e170f000801f8381c060f003e01f00000000f00f;
  defparam bm13.INIT_C = 256'h0000100804060200000000000000000000000e8783c1010000000787c3e10000;
  defparam bm13.INIT_D = 256'h000070381c0c0e00000038381c0e07000000381c0e0e070000001c1c0e870300;
  defparam bm13.INIT_E = 256'h0000c0e1707038000000c0e07038180000008040002010000000301008040200;
  defparam bm13.INIT_F = 256'h00000000000000000000808140603000000080c3e1e070000000c0c1e1703800;

  SB_RAM512x8 bm14 (
    .RDATA (data_int[14]),
    .RADDR (addr),
    .RCLK  (clk),
    .RCLKE (read_en[14]),
    .RE    (read_en[14]),
    .WADDR (9'h000),
    .WCLK  (1'b0),
    .WCLKE (1'b0),
    .WDATA (8'h00),
    .WE    (1'b0)
  );  
  defparam bm14.INIT_0 = 256'h00000000381c060000000000001c000000000000001c000000000000001c0000;
  defparam bm14.INIT_1 = 256'h000000f0807f80030000007030000607000000207008070200000000381c0e00;
  defparam bm14.INIT_2 = 256'h000000001e003e00000000807c801f00000000c0f9ffc700000000e0e1ffc301;
  defparam bm14.INIT_3 = 256'h0000fe003f00e0040000f8ff1f00f01e0000e0ff0700701e000000ff0f003808;
  defparam bm14.INIT_4 = 256'h00e001008003c0f900c00300c003c00100800f00f001c00100001f00fc00e000;
  defparam bm14.INIT_5 = 256'h00380000000ec00100700000000ec00100f00000000fc0f900e000008007c0fd;
  defparam bm14.INIT_6 = 256'h001f000000807f1e001c000000f8f71e0018000000fce30400380000003cc001;
  defparam bm14.INIT_7 = 256'h3c1c00000000e00ff81c00000000f807f01f00000000fc01c01f000000007e18;
  defparam bm14.INIT_8 = 256'h07380000000000700e380000000000780e1c00000000003c1c1c00000000001e;
  defparam bm14.INIT_9 = 256'h07e00000000000e007700000000000e007700000000000e007380000000000e0;
  defparam bm14.INIT_A = 256'h07001f00000000e007800700000000e007c00300000000e007e00100000000e0;
  defparam bm14.INIT_B = 256'h7800076f000e003c3c00e00f000000381c00f80f000000700e00fc00000000f0;
  defparam bm14.INIT_C = 256'h001ec761388e7300801f8761188ef303e01f0760000ef00ff0010760000e001f;
  defparam bm14.INIT_D = 256'h00000760000e00000000c761188e03000000c761388603000000c00138800300;
  defparam bm14.INIT_E = 256'h0000c261388403000000c001388003000000c761388e030000008761180e0300;
  defparam bm14.INIT_F = 256'h00000760000e000000000760000e000000000760000e00000000c761388e0300;

  SB_RAM512x8 bm15 (
    .RDATA (data_int[15]),
    .RADDR (addr),
    .RCLK  (clk),
    .RCLKE (read_en[15]),
    .RE    (read_en[15]),
    .WADDR (9'h000),
    .WCLK  (1'b0),
    .WCLKE (1'b0),
    .WDATA (8'h00),
    .WE    (1'b0)
  );  
  defparam bm15.INIT_0 = 256'h000000007338fc000000000073fc7f00000000001cfc1f00000000001cf80300;
  defparam bm15.INIT_1 = 256'h0000000000c0010f000000000ce08007000000001cf0c003000000003f78f001;
  defparam bm15.INIT_2 = 256'h000000007087037800000000f087033800000000c081013c00000000c0c1011e;
  defparam bm15.INIT_3 = 256'h0000fe003fc001e00000f8ffdf8003e00000e0ffc7810370000000fff0870370;
  defparam bm15.INIT_4 = 256'h00e0010080f300e000c00300c0e100e000800f00f0c101e000001f00fcc001e0;
  defparam bm15.INIT_5 = 256'h00380000001e00e000700000001e00e000f00000003f00e000e00000807f00c0;
  defparam bm15.INIT_6 = 256'h001f000000800f78001c000000f807700018000000fc037000380000003c00e0;
  defparam bm15.INIT_7 = 256'h3c1c00000000e00ff81c00000000f81ff01f00000000fc1dc01f000000001e38;
  defparam bm15.INIT_8 = 256'h07380000000000700e380000000000780e1c00000000003c1c1c00000000001e;
  defparam bm15.INIT_9 = 256'h07e00000000000e007700000000000e007700000000000e007380000000000e0;
  defparam bm15.INIT_A = 256'h07001f00000000e007800700000000e007c00300000000e007e00100000000e0;
  defparam bm15.INIT_B = 256'h7800076f000e003c3c00e00f000000381c00f80f000000700e00fc00000000f0;
  defparam bm15.INIT_C = 256'h001ec761388e7300801f8761188ef303e01f0760000ef00ff0010760000e001f;
  defparam bm15.INIT_D = 256'h00000760000e00000000c761188e03000000c761388603000000c00138800300;
  defparam bm15.INIT_E = 256'h0000c261388403000000c001388003000000c761388e030000008761180e0300;
  defparam bm15.INIT_F = 256'h00000760000e000000000760000e000000000760000e00000000c761388e0300; 

  SB_RAM512x8 bm16 (
    .RDATA (data_int[16]),
    .RADDR (addr),
    .RCLK  (clk),
    .RCLKE (read_en[16]),
    .RE    (read_en[16]),
    .WADDR (9'h000),
    .WCLK  (1'b0),
    .WCLKE (1'b0),
    .WDATA (8'h00),
    .WE    (1'b0)
  );  
  defparam bm16.INIT_0 = 256'h0000fcc13f0000000000f0ff0f0000000000c0ff030000000000001c00000000;
  defparam bm16.INIT_1 = 256'h00c00100c003000000c00700e001000000800f00f000000000003f007c000000;
  defparam bm16.INIT_2 = 256'h00380000000e000000700000000e000000f000000007000000e0010080070000;
  defparam bm16.INIT_3 = 256'h001e000000f80f00001c000000fc07000038000000fc010000380000001c0000;
  defparam bm16.INIT_4 = 256'h781c00000000f00ff01d00000000f803e01f00000000fc00c01f000000001e00;
  defparam bm16.INIT_5 = 256'h07380000000000700e180000000000381e1c00000000003c3c1c00000000001f;
  defparam bm16.INIT_6 = 256'h03e00000000000e007700000000000e007700000000000e007380000000000f0;
  defparam bm16.INIT_7 = 256'h07001f00000000e007800700000000e007c00300000000e007e00100000000c0;
  defparam bm16.INIT_8 = 256'h7800800f0000003c1c00f00f000000781e00f80f000000700e007e00000000e0;
  defparam bm16.INIT_9 = 256'h009f40000006f201c01f00000000f007e00f00000000e00ff80000000000001e;
  defparam bm16.INIT_A = 256'h0080c3011c0e0e0000c0e1001e0e070000c0e1000e0f070000e0600004870300;
  defparam bm16.INIT_B = 256'h00000e07f0783800000007037038180000000000380000000080c10038040600;
  defparam bm16.INIT_C = 256'h00000000fe03000000000c06ff61300000001c0ec0f1700000000e07e0703800;
  defparam bm16.INIT_D = 256'h0000e07038808703000070783c80c301000070381cc0c30100003018fe83c100;
  defparam bm16.INIT_E = 256'h000080c3c1011e0e000080c1e1000c0600000000f00000000000e07070008303;
  defparam bm16.INIT_F = 256'h0000000000000000000000878303381c0000008783033c1c000080c3c3031c0e;

  SB_RAM512x8 bm17 (
    .RDATA (data_int[17]),
    .RADDR (addr),
    .RCLK  (clk),
    .RCLKE (read_en[17]),
    .RE    (read_en[17]),
    .WADDR (9'h000),
    .WCLK  (1'b0),
    .WCLKE (1'b0),
    .WDATA (8'h00),
    .WE    (1'b0)
  );  
  defparam bm17.INIT_0 = 256'h00003e007e0000000000fcf71f0000000000f0ff07000000000080ff01000000;
  defparam bm17.INIT_1 = 256'h00e001008007000000c00300c003000000800700e001000000001f00f8000000;
  defparam bm17.INIT_2 = 256'h00380000001e000000780000000e000000700000000e000000f0000000070000;
  defparam bm17.INIT_3 = 256'h801f000000001f00001c000000f80f00001c000000fc03000038000000fc0000;
  defparam bm17.INIT_4 = 256'h3c1c00000000801f781c00000000f007f01d00000000f803e01f000000007c00;
  defparam bm17.INIT_5 = 256'h07380000000000700f380000000000700e1c0000000000381c1c00000000003e;
  defparam bm17.INIT_6 = 256'h07e00100000000e007f00000000000e007700000000000e007780000000000e0;
  defparam bm17.INIT_7 = 256'h0e003e00000000e007000f00000000e007800700000000e007c00300000000e0;
  defparam bm17.INIT_8 = 256'hf80000000000001e3c00c00f0000003c1c00f00f000000780e00fc0300000070;
  defparam bm17.INIT_9 = 256'h00f8ffffffff1f0080ffffffffffff01c0ffffffffffff07f00700000000c00f;
  defparam bm17.INIT_A = 256'h0080ff0000ff01000000dd0000bb000000001c00003800000000000000000000;
  defparam bm17.INIT_B = 256'h0080fff81fff01000080ff9009ff010000007f8001fe00000080ff0000ff0100;
  defparam bm17.INIT_C = 256'h00001cf81f380000000000f81f00000000001ce00738000000009df81fb90000;
  defparam bm17.INIT_D = 256'h00007f8001fe00000080ff0000ff01000080ff8001ff010000001c9009380000;
  defparam bm17.INIT_E = 256'h00001cf00f3800000080ddf81fbb01000080fff00fff01000080ff8001ff0100;
  defparam bm17.INIT_F = 256'h0000008001000000000000b00d000000000000f81f000000000000f00f000000; 

  SB_RAM512x8 bm18 (
    .RDATA (data_int[18]),
    .RADDR (addr),
    .RCLK  (clk),
    .RCLKE (read_en[18]),
    .RE    (read_en[18]),
    .WADDR (9'h000),
    .WCLK  (1'b0),
    .WCLKE (1'b0),
    .WDATA (8'h00),
    .WE    (1'b0)
  );  
  defparam bm18.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam bm18.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam bm18.INIT_2 = 256'h7ffe9ffff3fffc7ffc3fffc7fff13ffcf80ffc837fe01ff8e007f8003ec00fe0;
  defparam bm18.INIT_3 = 256'h000000000000000002c00010000480000ff003fe801fe0071ffc07ffc17ff81f;
  defparam bm18.INIT_4 = 256'hf00ffc017fc00ff0c00370001c0003c000000000000000000000000000000000;
  defparam bm18.INIT_5 = 256'h0ff807fec03ff00f3ffc0fffe37ff83ffeffffefffff7f7ffc1ffe87fff03ff8;
  defparam bm18.INIT_6 = 256'h00000000000000000000000000000000000000000000000007e00178000fc003;
  defparam bm18.INIT_7 = 256'hfc3fffc7fff97ffef80ffc83ffe01ff8e007f8013ec00fe00000000000000000;
  defparam bm18.INIT_8 = 256'h000000000000000007f0037c801fe0071ff807ffc13ff81f7ffe9fffe3fffc3f;
  defparam bm18.INIT_9 = 256'hc003f0001e8007e0000000000000000000000000000000000000000000000000;
  defparam bm18.INIT_A = 256'h1ffc0fffe17ff83ffeffdffff7ffff7ffc1ffec7fff03ffcf00ffc017fe01ff0;
  defparam bm18.INIT_B = 256'h0000000000000000000000000000000003c00038000ec0030ff003fe803ff00f;
  defparam bm18.INIT_C = 256'hf81ffe83ffe01ff8f007f8013fc00ff080012000080003400000000000000000;
  defparam bm18.INIT_D = 256'h07f0037c001fe0070ff807fec13ff01f3ffc8fffe3fffc3ffe3fffeffff97ffe;
  defparam bm18.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  defparam bm18.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
  
endmodule  